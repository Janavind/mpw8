magic
tech sky130A
magscale 1 2
timestamp 1672275371
<< viali >>
rect 3433 57545 3467 57579
rect 5273 57545 5307 57579
rect 10793 57545 10827 57579
rect 12173 57545 12207 57579
rect 13553 57545 13587 57579
rect 14933 57545 14967 57579
rect 16957 57545 16991 57579
rect 17693 57545 17727 57579
rect 19533 57545 19567 57579
rect 20453 57545 20487 57579
rect 22293 57545 22327 57579
rect 26065 57545 26099 57579
rect 27445 57545 27479 57579
rect 28733 57545 28767 57579
rect 39405 57545 39439 57579
rect 54033 57545 54067 57579
rect 55597 57545 55631 57579
rect 4077 57477 4111 57511
rect 31677 57477 31711 57511
rect 33977 57477 34011 57511
rect 45845 57477 45879 57511
rect 53021 57477 53055 57511
rect 5457 57409 5491 57443
rect 7297 57409 7331 57443
rect 7757 57409 7791 57443
rect 8585 57409 8619 57443
rect 9321 57409 9355 57443
rect 10057 57409 10091 57443
rect 10977 57409 11011 57443
rect 12357 57409 12391 57443
rect 12817 57409 12851 57443
rect 13737 57409 13771 57443
rect 15117 57409 15151 57443
rect 15761 57409 15795 57443
rect 17141 57409 17175 57443
rect 17877 57409 17911 57443
rect 18521 57409 18555 57443
rect 19717 57409 19751 57443
rect 20637 57409 20671 57443
rect 22477 57409 22511 57443
rect 23213 57409 23247 57443
rect 23673 57409 23707 57443
rect 23857 57409 23891 57443
rect 24777 57409 24811 57443
rect 25881 57409 25915 57443
rect 27261 57409 27295 57443
rect 27997 57409 28031 57443
rect 28181 57409 28215 57443
rect 28917 57409 28951 57443
rect 30205 57409 30239 57443
rect 30849 57409 30883 57443
rect 33793 57409 33827 57443
rect 34069 57409 34103 57443
rect 35357 57409 35391 57443
rect 35541 57409 35575 57443
rect 36001 57409 36035 57443
rect 37473 57409 37507 57443
rect 40049 57409 40083 57443
rect 40325 57409 40359 57443
rect 41521 57409 41555 57443
rect 43729 57409 43763 57443
rect 44373 57409 44407 57443
rect 44649 57409 44683 57443
rect 49065 57409 49099 57443
rect 50353 57409 50387 57443
rect 50629 57409 50663 57443
rect 51641 57409 51675 57443
rect 54217 57409 54251 57443
rect 54677 57409 54711 57443
rect 55781 57409 55815 57443
rect 56885 57409 56919 57443
rect 6009 57341 6043 57375
rect 24961 57341 24995 57375
rect 31493 57341 31527 57375
rect 32321 57341 32355 57375
rect 32597 57341 32631 57375
rect 36277 57341 36311 57375
rect 37749 57341 37783 57375
rect 41797 57341 41831 57375
rect 43453 57341 43487 57375
rect 44557 57341 44591 57375
rect 47777 57341 47811 57375
rect 56241 57341 56275 57375
rect 4261 57273 4295 57307
rect 23029 57273 23063 57307
rect 24593 57273 24627 57307
rect 30389 57273 30423 57307
rect 35173 57273 35207 57307
rect 41705 57273 41739 57307
rect 49709 57273 49743 57307
rect 21465 57205 21499 57239
rect 24041 57205 24075 57239
rect 28181 57205 28215 57239
rect 33609 57205 33643 57239
rect 38761 57205 38795 57239
rect 41337 57205 41371 57239
rect 44189 57205 44223 57239
rect 45753 57205 45787 57239
rect 46397 57205 46431 57239
rect 47041 57205 47075 57239
rect 48007 57205 48041 57239
rect 51825 57205 51859 57239
rect 53113 57205 53147 57239
rect 4721 57001 4755 57035
rect 5917 57001 5951 57035
rect 6561 57001 6595 57035
rect 11621 57001 11655 57035
rect 14381 57001 14415 57035
rect 17141 57001 17175 57035
rect 19901 57001 19935 57035
rect 21097 57001 21131 57035
rect 21833 57001 21867 57035
rect 23489 57001 23523 57035
rect 24041 57001 24075 57035
rect 27261 57001 27295 57035
rect 27721 57001 27755 57035
rect 31309 57001 31343 57035
rect 41061 57001 41095 57035
rect 41613 57001 41647 57035
rect 42901 57001 42935 57035
rect 47777 57001 47811 57035
rect 50353 57001 50387 57035
rect 50997 57001 51031 57035
rect 51641 57001 51675 57035
rect 52285 57001 52319 57035
rect 53021 57001 53055 57035
rect 53665 57001 53699 57035
rect 54309 57001 54343 57035
rect 56149 57001 56183 57035
rect 11161 56933 11195 56967
rect 22937 56933 22971 56967
rect 28549 56933 28583 56967
rect 28825 56933 28859 56967
rect 31769 56933 31803 56967
rect 33241 56933 33275 56967
rect 36369 56933 36403 56967
rect 39313 56933 39347 56967
rect 43453 56933 43487 56967
rect 47133 56933 47167 56967
rect 23397 56865 23431 56899
rect 25053 56865 25087 56899
rect 29009 56865 29043 56899
rect 29745 56865 29779 56899
rect 30205 56865 30239 56899
rect 35081 56865 35115 56899
rect 35265 56865 35299 56899
rect 38025 56865 38059 56899
rect 38209 56865 38243 56899
rect 40325 56865 40359 56899
rect 40509 56865 40543 56899
rect 41705 56865 41739 56899
rect 43361 56865 43395 56899
rect 46489 56865 46523 56899
rect 48421 56865 48455 56899
rect 49709 56865 49743 56899
rect 22017 56797 22051 56831
rect 23903 56797 23937 56831
rect 25145 56797 25179 56831
rect 25516 56797 25550 56831
rect 26617 56797 26651 56831
rect 26801 56797 26835 56831
rect 27445 56797 27479 56831
rect 27537 56797 27571 56831
rect 27813 56797 27847 56831
rect 28733 56797 28767 56831
rect 28917 56797 28951 56831
rect 29193 56797 29227 56831
rect 29929 56797 29963 56831
rect 30113 56797 30147 56831
rect 30297 56797 30331 56831
rect 30481 56797 30515 56831
rect 31894 56797 31928 56831
rect 32321 56797 32355 56831
rect 32413 56797 32447 56831
rect 33057 56797 33091 56831
rect 33333 56797 33367 56831
rect 33977 56797 34011 56831
rect 34161 56797 34195 56831
rect 34253 56797 34287 56831
rect 35449 56797 35483 56831
rect 35633 56797 35667 56831
rect 36277 56797 36311 56831
rect 36553 56797 36587 56831
rect 36737 56797 36771 56831
rect 37013 56797 37047 56831
rect 38301 56797 38335 56831
rect 38393 56797 38427 56831
rect 38485 56797 38519 56831
rect 39037 56797 39071 56831
rect 40233 56797 40267 56831
rect 40417 56797 40451 56831
rect 41186 56797 41220 56831
rect 42165 56797 42199 56831
rect 43545 56797 43579 56831
rect 43913 56797 43947 56831
rect 44189 56797 44223 56831
rect 45201 56797 45235 56831
rect 46029 56797 46063 56831
rect 48697 56797 48731 56831
rect 55505 56797 55539 56831
rect 26709 56729 26743 56763
rect 33793 56729 33827 56763
rect 39313 56729 39347 56763
rect 23857 56661 23891 56695
rect 25513 56661 25547 56695
rect 25697 56661 25731 56695
rect 31953 56661 31987 56695
rect 32873 56661 32907 56695
rect 39129 56661 39163 56695
rect 40049 56661 40083 56695
rect 41245 56661 41279 56695
rect 45845 56661 45879 56695
rect 23397 56457 23431 56491
rect 27629 56457 27663 56491
rect 28273 56457 28307 56491
rect 29101 56457 29135 56491
rect 30849 56457 30883 56491
rect 32597 56457 32631 56491
rect 43729 56457 43763 56491
rect 50169 56457 50203 56491
rect 51457 56457 51491 56491
rect 53021 56457 53055 56491
rect 36461 56389 36495 56423
rect 36829 56389 36863 56423
rect 40325 56389 40359 56423
rect 40417 56389 40451 56423
rect 44097 56389 44131 56423
rect 22661 56321 22695 56355
rect 23581 56321 23615 56355
rect 24041 56321 24075 56355
rect 25421 56321 25455 56355
rect 26249 56321 26283 56355
rect 26433 56321 26467 56355
rect 27261 56321 27295 56355
rect 27688 56321 27722 56355
rect 28457 56321 28491 56355
rect 28641 56321 28675 56355
rect 29101 56321 29135 56355
rect 29377 56321 29411 56355
rect 30021 56321 30055 56355
rect 31217 56321 31251 56355
rect 31309 56321 31343 56355
rect 32689 56321 32723 56355
rect 33333 56321 33367 56355
rect 33425 56321 33459 56355
rect 33609 56321 33643 56355
rect 33701 56321 33735 56355
rect 34161 56321 34195 56355
rect 34345 56321 34379 56355
rect 34621 56321 34655 56355
rect 35724 56321 35758 56355
rect 35817 56321 35851 56355
rect 36645 56321 36679 56355
rect 36921 56321 36955 56355
rect 38853 56321 38887 56355
rect 40187 56321 40221 56355
rect 40509 56321 40543 56355
rect 41613 56321 41647 56355
rect 42625 56321 42659 56355
rect 42809 56321 42843 56355
rect 42901 56321 42935 56355
rect 43085 56321 43119 56355
rect 43177 56321 43211 56355
rect 43637 56321 43671 56355
rect 43913 56321 43947 56355
rect 44925 56321 44959 56355
rect 45783 56321 45817 56355
rect 45937 56321 45971 56355
rect 47041 56321 47075 56355
rect 47961 56321 47995 56355
rect 48881 56321 48915 56355
rect 49525 56321 49559 56355
rect 24317 56253 24351 56287
rect 25237 56253 25271 56287
rect 26617 56253 26651 56287
rect 27169 56253 27203 56287
rect 29193 56253 29227 56287
rect 31033 56253 31067 56287
rect 31125 56253 31159 56287
rect 38209 56253 38243 56287
rect 38669 56253 38703 56287
rect 39037 56253 39071 56287
rect 40049 56253 40083 56287
rect 40693 56253 40727 56287
rect 41889 56253 41923 56287
rect 44833 56253 44867 56287
rect 27813 56185 27847 56219
rect 37933 56185 37967 56219
rect 44557 56185 44591 56219
rect 46397 56185 46431 56219
rect 25605 56117 25639 56151
rect 33149 56117 33183 56151
rect 34529 56117 34563 56151
rect 35633 56117 35667 56151
rect 37749 56117 37783 56151
rect 39589 56117 39623 56151
rect 41429 56117 41463 56151
rect 41797 56117 41831 56151
rect 45753 56117 45787 56151
rect 23857 55913 23891 55947
rect 24685 55913 24719 55947
rect 27997 55913 28031 55947
rect 31585 55913 31619 55947
rect 34345 55913 34379 55947
rect 35909 55913 35943 55947
rect 37013 55913 37047 55947
rect 37657 55913 37691 55947
rect 39037 55913 39071 55947
rect 40049 55913 40083 55947
rect 41613 55913 41647 55947
rect 42625 55913 42659 55947
rect 42993 55913 43027 55947
rect 43453 55913 43487 55947
rect 46857 55913 46891 55947
rect 32965 55845 32999 55879
rect 34897 55845 34931 55879
rect 40877 55845 40911 55879
rect 44373 55845 44407 55879
rect 45477 55845 45511 55879
rect 45569 55845 45603 55879
rect 23397 55777 23431 55811
rect 25697 55777 25731 55811
rect 26249 55777 26283 55811
rect 26709 55777 26743 55811
rect 28641 55777 28675 55811
rect 28733 55777 28767 55811
rect 29929 55777 29963 55811
rect 33425 55777 33459 55811
rect 35173 55777 35207 55811
rect 36829 55777 36863 55811
rect 24041 55709 24075 55743
rect 24869 55709 24903 55743
rect 25329 55709 25363 55743
rect 25513 55709 25547 55743
rect 26893 55709 26927 55743
rect 27721 55709 27755 55743
rect 27997 55709 28031 55743
rect 28549 55709 28583 55743
rect 28825 55709 28859 55743
rect 30941 55709 30975 55743
rect 31217 55709 31251 55743
rect 31401 55709 31435 55743
rect 32229 55709 32263 55743
rect 32505 55709 32539 55743
rect 33149 55709 33183 55743
rect 33333 55709 33367 55743
rect 34069 55709 34103 55743
rect 34161 55709 34195 55743
rect 34345 55709 34379 55743
rect 35265 55709 35299 55743
rect 36737 55709 36771 55743
rect 38117 55709 38151 55743
rect 38301 55709 38335 55743
rect 38577 55709 38611 55743
rect 42533 55709 42567 55743
rect 42809 55709 42843 55743
rect 44097 55709 44131 55743
rect 44373 55709 44407 55743
rect 45201 55709 45235 55743
rect 45385 55709 45419 55743
rect 45661 55709 45695 55743
rect 27813 55641 27847 55675
rect 30113 55641 30147 55675
rect 30297 55641 30331 55675
rect 31079 55641 31113 55675
rect 31309 55641 31343 55675
rect 32045 55641 32079 55675
rect 32413 55641 32447 55675
rect 39221 55641 39255 55675
rect 39405 55641 39439 55675
rect 40233 55641 40267 55675
rect 40417 55641 40451 55675
rect 41797 55641 41831 55675
rect 41981 55641 42015 55675
rect 27077 55573 27111 55607
rect 29009 55573 29043 55607
rect 38485 55573 38519 55607
rect 44189 55573 44223 55607
rect 46213 55573 46247 55607
rect 23949 55369 23983 55403
rect 25697 55369 25731 55403
rect 26433 55369 26467 55403
rect 27353 55369 27387 55403
rect 27997 55369 28031 55403
rect 30941 55369 30975 55403
rect 32321 55369 32355 55403
rect 34437 55369 34471 55403
rect 35081 55369 35115 55403
rect 40147 55369 40181 55403
rect 44281 55369 44315 55403
rect 46213 55369 46247 55403
rect 24501 55301 24535 55335
rect 25053 55301 25087 55335
rect 29101 55301 29135 55335
rect 39221 55301 39255 55335
rect 45753 55301 45787 55335
rect 25513 55233 25547 55267
rect 26617 55233 26651 55267
rect 27169 55233 27203 55267
rect 27813 55233 27847 55267
rect 29285 55233 29319 55267
rect 29377 55233 29411 55267
rect 30021 55233 30055 55267
rect 30205 55233 30239 55267
rect 31125 55233 31159 55267
rect 31309 55233 31343 55267
rect 32505 55233 32539 55267
rect 32689 55233 32723 55267
rect 34621 55233 34655 55267
rect 35265 55233 35299 55267
rect 35541 55233 35575 55267
rect 38209 55233 38243 55267
rect 38301 55233 38335 55267
rect 38485 55233 38519 55267
rect 38577 55233 38611 55267
rect 39405 55233 39439 55267
rect 39589 55233 39623 55267
rect 40049 55233 40083 55267
rect 40233 55233 40267 55267
rect 40325 55233 40359 55267
rect 41797 55233 41831 55267
rect 42901 55233 42935 55267
rect 42993 55233 43027 55267
rect 43121 55233 43155 55267
rect 43637 55233 43671 55267
rect 44465 55233 44499 55267
rect 44925 55233 44959 55267
rect 28641 55165 28675 55199
rect 33793 55165 33827 55199
rect 36093 55165 36127 55199
rect 36737 55165 36771 55199
rect 37473 55165 37507 55199
rect 38761 55165 38795 55199
rect 40785 55165 40819 55199
rect 33149 55097 33183 55131
rect 35357 55097 35391 55131
rect 35449 55097 35483 55131
rect 29101 55029 29135 55063
rect 29837 55029 29871 55063
rect 41337 55029 41371 55063
rect 41705 55029 41739 55063
rect 42717 55029 42751 55063
rect 25145 54825 25179 54859
rect 25789 54825 25823 54859
rect 26525 54825 26559 54859
rect 27905 54825 27939 54859
rect 30297 54825 30331 54859
rect 30849 54825 30883 54859
rect 31953 54825 31987 54859
rect 32873 54825 32907 54859
rect 33609 54825 33643 54859
rect 33793 54825 33827 54859
rect 34897 54825 34931 54859
rect 35633 54825 35667 54859
rect 36185 54825 36219 54859
rect 37289 54825 37323 54859
rect 38117 54825 38151 54859
rect 39497 54825 39531 54859
rect 40877 54825 40911 54859
rect 41705 54825 41739 54859
rect 28457 54757 28491 54791
rect 36737 54757 36771 54791
rect 40049 54757 40083 54791
rect 43729 54757 43763 54791
rect 28825 54689 28859 54723
rect 39221 54689 39255 54723
rect 41245 54689 41279 54723
rect 42809 54689 42843 54723
rect 42901 54689 42935 54723
rect 43269 54689 43303 54723
rect 44189 54689 44223 54723
rect 26985 54621 27019 54655
rect 29745 54621 29779 54655
rect 29837 54621 29871 54655
rect 30021 54621 30055 54655
rect 30113 54621 30147 54655
rect 30849 54621 30883 54655
rect 31033 54621 31067 54655
rect 31125 54621 31159 54655
rect 31769 54621 31803 54655
rect 33149 54621 33183 54655
rect 38301 54621 38335 54655
rect 38485 54621 38519 54655
rect 39129 54621 39163 54655
rect 40785 54621 40819 54655
rect 41889 54621 41923 54655
rect 42165 54621 42199 54655
rect 44097 54621 44131 54655
rect 27077 54553 27111 54587
rect 33761 54553 33795 54587
rect 33977 54553 34011 54587
rect 28365 54485 28399 54519
rect 32229 54485 32263 54519
rect 32689 54485 32723 54519
rect 42073 54485 42107 54519
rect 42625 54485 42659 54519
rect 26525 54281 26559 54315
rect 27169 54281 27203 54315
rect 27813 54281 27847 54315
rect 28273 54281 28307 54315
rect 29377 54281 29411 54315
rect 31217 54281 31251 54315
rect 32873 54281 32907 54315
rect 34345 54281 34379 54315
rect 36461 54281 36495 54315
rect 37473 54281 37507 54315
rect 39129 54281 39163 54315
rect 40509 54281 40543 54315
rect 41521 54281 41555 54315
rect 41981 54281 42015 54315
rect 42717 54281 42751 54315
rect 44189 54281 44223 54315
rect 29561 54213 29595 54247
rect 35909 54213 35943 54247
rect 43085 54213 43119 54247
rect 28641 54145 28675 54179
rect 29745 54145 29779 54179
rect 30389 54145 30423 54179
rect 32505 54145 32539 54179
rect 33885 54145 33919 54179
rect 35173 54145 35207 54179
rect 39221 54145 39255 54179
rect 39681 54145 39715 54179
rect 40325 54145 40359 54179
rect 41153 54145 41187 54179
rect 42625 54145 42659 54179
rect 42901 54145 42935 54179
rect 43821 54145 43855 54179
rect 44005 54145 44039 54179
rect 28549 54077 28583 54111
rect 30481 54077 30515 54111
rect 30757 54077 30791 54111
rect 32413 54077 32447 54111
rect 33977 54077 34011 54111
rect 35081 54077 35115 54111
rect 41245 54077 41279 54111
rect 43729 54077 43763 54111
rect 33701 53941 33735 53975
rect 34897 53941 34931 53975
rect 27905 53737 27939 53771
rect 29929 53737 29963 53771
rect 30757 53737 30791 53771
rect 31953 53737 31987 53771
rect 32873 53737 32907 53771
rect 33885 53737 33919 53771
rect 34897 53737 34931 53771
rect 35265 53737 35299 53771
rect 35909 53737 35943 53771
rect 40233 53737 40267 53771
rect 42073 53737 42107 53771
rect 42257 53737 42291 53771
rect 26985 53669 27019 53703
rect 29193 53669 29227 53703
rect 31401 53669 31435 53703
rect 39405 53669 39439 53703
rect 40785 53669 40819 53703
rect 41337 53669 41371 53703
rect 30297 53601 30331 53635
rect 35357 53601 35391 53635
rect 30113 53533 30147 53567
rect 32137 53533 32171 53567
rect 32413 53533 32447 53567
rect 33057 53533 33091 53567
rect 33333 53533 33367 53567
rect 34069 53533 34103 53567
rect 34171 53533 34205 53567
rect 34289 53533 34323 53567
rect 35081 53533 35115 53567
rect 32321 53465 32355 53499
rect 33241 53465 33275 53499
rect 42441 53465 42475 53499
rect 42241 53397 42275 53431
rect 30481 53193 30515 53227
rect 31493 53193 31527 53227
rect 32781 53193 32815 53227
rect 33333 53193 33367 53227
rect 33885 53193 33919 53227
rect 34437 53193 34471 53227
rect 39865 53193 39899 53227
rect 32137 52649 32171 52683
rect 34345 52037 34379 52071
rect 34161 51901 34195 51935
rect 35725 51901 35759 51935
rect 34161 51561 34195 51595
rect 29561 8585 29595 8619
rect 30481 8449 30515 8483
rect 30573 8313 30607 8347
rect 27813 7837 27847 7871
rect 29009 7837 29043 7871
rect 29929 7837 29963 7871
rect 30481 7837 30515 7871
rect 31309 7837 31343 7871
rect 27905 7701 27939 7735
rect 29101 7701 29135 7735
rect 29837 7701 29871 7735
rect 31217 7701 31251 7735
rect 29561 7429 29595 7463
rect 28917 7293 28951 7327
rect 29377 7293 29411 7327
rect 30757 7293 30791 7327
rect 27353 7157 27387 7191
rect 27997 7157 28031 7191
rect 27353 6817 27387 6851
rect 27537 6817 27571 6851
rect 28089 6817 28123 6851
rect 31125 6817 31159 6851
rect 31677 6817 31711 6851
rect 24869 6749 24903 6783
rect 25513 6749 25547 6783
rect 26709 6749 26743 6783
rect 29745 6749 29779 6783
rect 30941 6749 30975 6783
rect 33793 6749 33827 6783
rect 30021 6681 30055 6715
rect 25421 6613 25455 6647
rect 26249 6613 26283 6647
rect 26801 6613 26835 6647
rect 32965 6409 32999 6443
rect 29377 6341 29411 6375
rect 26433 6273 26467 6307
rect 27261 6273 27295 6307
rect 31493 6273 31527 6307
rect 35357 6273 35391 6307
rect 27445 6205 27479 6239
rect 29193 6205 29227 6239
rect 29745 6205 29779 6239
rect 33885 6205 33919 6239
rect 35173 6205 35207 6239
rect 25421 6069 25455 6103
rect 26525 6069 26559 6103
rect 28733 6069 28767 6103
rect 32505 6069 32539 6103
rect 35633 5865 35667 5899
rect 25053 5729 25087 5763
rect 25237 5729 25271 5763
rect 25973 5729 26007 5763
rect 27353 5729 27387 5763
rect 27537 5729 27571 5763
rect 27813 5729 27847 5763
rect 30481 5729 30515 5763
rect 30665 5729 30699 5763
rect 31401 5729 31435 5763
rect 30021 5661 30055 5695
rect 32781 5661 32815 5695
rect 33057 5661 33091 5695
rect 33701 5661 33735 5695
rect 34897 5661 34931 5695
rect 35725 5661 35759 5695
rect 36369 5661 36403 5695
rect 33793 5525 33827 5559
rect 36277 5525 36311 5559
rect 27353 5253 27387 5287
rect 33977 5253 34011 5287
rect 36277 5253 36311 5287
rect 29469 5185 29503 5219
rect 34161 5185 34195 5219
rect 26617 5117 26651 5151
rect 27169 5117 27203 5151
rect 27721 5117 27755 5151
rect 29653 5117 29687 5151
rect 30389 5117 30423 5151
rect 32505 5117 32539 5151
rect 34713 5117 34747 5151
rect 36461 5117 36495 5151
rect 23765 4981 23799 5015
rect 24685 4981 24719 5015
rect 25329 4981 25363 5015
rect 25973 4981 26007 5015
rect 29193 4777 29227 4811
rect 36369 4777 36403 4811
rect 23397 4709 23431 4743
rect 25513 4709 25547 4743
rect 26617 4641 26651 4675
rect 27629 4641 27663 4675
rect 29929 4641 29963 4675
rect 30573 4641 30607 4675
rect 32689 4641 32723 4675
rect 34069 4641 34103 4675
rect 21557 4573 21591 4607
rect 22385 4573 22419 4607
rect 23857 4573 23891 4607
rect 24685 4573 24719 4607
rect 26157 4573 26191 4607
rect 35081 4573 35115 4607
rect 35541 4573 35575 4607
rect 36829 4573 36863 4607
rect 23949 4505 23983 4539
rect 26801 4505 26835 4539
rect 30113 4505 30147 4539
rect 33885 4505 33919 4539
rect 34989 4505 35023 4539
rect 24777 4437 24811 4471
rect 23489 4097 23523 4131
rect 24777 4097 24811 4131
rect 27629 4097 27663 4131
rect 29929 4097 29963 4131
rect 34989 4097 35023 4131
rect 35817 4097 35851 4131
rect 23581 4029 23615 4063
rect 24961 4029 24995 4063
rect 26433 4029 26467 4063
rect 27813 4029 27847 4063
rect 28365 4029 28399 4063
rect 30113 4029 30147 4063
rect 30849 4029 30883 4063
rect 33057 4029 33091 4063
rect 34345 4029 34379 4063
rect 34529 4029 34563 4063
rect 37473 4029 37507 4063
rect 22385 3961 22419 3995
rect 35725 3961 35759 3995
rect 38117 3961 38151 3995
rect 17417 3893 17451 3927
rect 19625 3893 19659 3927
rect 20453 3893 20487 3927
rect 21465 3893 21499 3927
rect 23029 3893 23063 3927
rect 24317 3893 24351 3927
rect 35081 3893 35115 3927
rect 36277 3893 36311 3927
rect 38761 3893 38795 3927
rect 39497 3893 39531 3927
rect 22109 3689 22143 3723
rect 29837 3689 29871 3723
rect 30481 3689 30515 3723
rect 37841 3689 37875 3723
rect 21465 3621 21499 3655
rect 38485 3621 38519 3655
rect 40049 3621 40083 3655
rect 41981 3621 42015 3655
rect 45845 3621 45879 3655
rect 47777 3621 47811 3655
rect 20821 3553 20855 3587
rect 22753 3553 22787 3587
rect 25237 3553 25271 3587
rect 26709 3553 26743 3587
rect 27353 3553 27387 3587
rect 28917 3553 28951 3587
rect 32229 3553 32263 3587
rect 34897 3553 34931 3587
rect 36737 3553 36771 3587
rect 40693 3553 40727 3587
rect 42625 3553 42659 3587
rect 43913 3553 43947 3587
rect 9137 3485 9171 3519
rect 10057 3485 10091 3519
rect 10885 3485 10919 3519
rect 11713 3485 11747 3519
rect 12541 3485 12575 3519
rect 13369 3485 13403 3519
rect 14289 3485 14323 3519
rect 15025 3485 15059 3519
rect 15853 3485 15887 3519
rect 16681 3485 16715 3519
rect 17601 3485 17635 3519
rect 18245 3485 18279 3519
rect 18889 3485 18923 3519
rect 20177 3485 20211 3519
rect 23397 3485 23431 3519
rect 23857 3485 23891 3519
rect 25053 3485 25087 3519
rect 29929 3485 29963 3519
rect 30573 3485 30607 3519
rect 33425 3485 33459 3519
rect 33885 3485 33919 3519
rect 37381 3485 37415 3519
rect 39129 3485 39163 3519
rect 41337 3485 41371 3519
rect 43269 3485 43303 3519
rect 45201 3485 45235 3519
rect 46489 3485 46523 3519
rect 47133 3485 47167 3519
rect 48421 3485 48455 3519
rect 49157 3485 49191 3519
rect 50537 3485 50571 3519
rect 51181 3485 51215 3519
rect 51825 3485 51859 3519
rect 27537 3417 27571 3451
rect 33241 3417 33275 3451
rect 36553 3417 36587 3451
rect 37289 3417 37323 3451
rect 23949 3349 23983 3383
rect 24225 3077 24259 3111
rect 33977 3077 34011 3111
rect 36277 3077 36311 3111
rect 38209 3077 38243 3111
rect 20821 3009 20855 3043
rect 21465 3009 21499 3043
rect 22385 3009 22419 3043
rect 22845 3009 22879 3043
rect 24133 3009 24167 3043
rect 24777 3009 24811 3043
rect 34161 3009 34195 3043
rect 37657 3009 37691 3043
rect 38117 3009 38151 3043
rect 39405 3009 39439 3043
rect 43913 3009 43947 3043
rect 13737 2941 13771 2975
rect 15669 2941 15703 2975
rect 19533 2941 19567 2975
rect 24961 2941 24995 2975
rect 26617 2941 26651 2975
rect 27629 2941 27663 2975
rect 27813 2941 27847 2975
rect 29193 2941 29227 2975
rect 29929 2941 29963 2975
rect 30113 2941 30147 2975
rect 31125 2941 31159 2975
rect 32321 2941 32355 2975
rect 34621 2941 34655 2975
rect 36461 2941 36495 2975
rect 38761 2941 38795 2975
rect 40693 2941 40727 2975
rect 42625 2941 42659 2975
rect 44557 2941 44591 2975
rect 45845 2941 45879 2975
rect 49709 2941 49743 2975
rect 18889 2873 18923 2907
rect 20177 2873 20211 2907
rect 23673 2873 23707 2907
rect 41337 2873 41371 2907
rect 46489 2873 46523 2907
rect 48421 2873 48455 2907
rect 50353 2873 50387 2907
rect 51641 2873 51675 2907
rect 8309 2805 8343 2839
rect 9229 2805 9263 2839
rect 9873 2805 9907 2839
rect 10517 2805 10551 2839
rect 11161 2805 11195 2839
rect 12449 2805 12483 2839
rect 13093 2805 13127 2839
rect 14381 2805 14415 2839
rect 15025 2805 15059 2839
rect 16313 2805 16347 2839
rect 17601 2805 17635 2839
rect 18245 2805 18279 2839
rect 22937 2805 22971 2839
rect 37565 2805 37599 2839
rect 40049 2805 40083 2839
rect 43269 2805 43303 2839
rect 45201 2805 45235 2839
rect 47777 2805 47811 2839
rect 49065 2805 49099 2839
rect 50997 2805 51031 2839
rect 52929 2805 52963 2839
rect 23305 2601 23339 2635
rect 23949 2601 23983 2635
rect 34989 2601 35023 2635
rect 37473 2601 37507 2635
rect 38761 2601 38795 2635
rect 40049 2601 40083 2635
rect 7941 2533 7975 2567
rect 9873 2533 9907 2567
rect 13737 2533 13771 2567
rect 15669 2533 15703 2567
rect 17601 2533 17635 2567
rect 22661 2533 22695 2567
rect 25329 2533 25363 2567
rect 35541 2533 35575 2567
rect 43913 2533 43947 2567
rect 46489 2533 46523 2567
rect 50353 2533 50387 2567
rect 53573 2533 53607 2567
rect 13093 2465 13127 2499
rect 16313 2465 16347 2499
rect 18245 2465 18279 2499
rect 20177 2465 20211 2499
rect 27353 2465 27387 2499
rect 27537 2465 27571 2499
rect 28549 2465 28583 2499
rect 29745 2465 29779 2499
rect 30205 2465 30239 2499
rect 33333 2465 33367 2499
rect 34345 2465 34379 2499
rect 40693 2465 40727 2499
rect 43269 2465 43303 2499
rect 45201 2465 45235 2499
rect 48421 2465 48455 2499
rect 50997 2465 51031 2499
rect 54217 2465 54251 2499
rect 7297 2397 7331 2431
rect 8585 2397 8619 2431
rect 10517 2397 10551 2431
rect 11161 2397 11195 2431
rect 12449 2397 12483 2431
rect 15025 2397 15059 2431
rect 18889 2397 18923 2431
rect 20821 2397 20855 2431
rect 21465 2397 21499 2431
rect 22753 2397 22787 2431
rect 23213 2397 23247 2431
rect 24041 2397 24075 2431
rect 25789 2397 25823 2431
rect 26617 2397 26651 2431
rect 35081 2397 35115 2431
rect 36369 2397 36403 2431
rect 38117 2397 38151 2431
rect 41337 2397 41371 2431
rect 42625 2397 42659 2431
rect 45845 2397 45879 2431
rect 47777 2397 47811 2431
rect 49065 2397 49099 2431
rect 51641 2397 51675 2431
rect 52929 2397 52963 2431
rect 29929 2329 29963 2363
rect 34161 2329 34195 2363
rect 36277 2329 36311 2363
rect 25881 2261 25915 2295
<< metal1 >>
rect 21358 57876 21364 57928
rect 21416 57916 21422 57928
rect 27430 57916 27436 57928
rect 21416 57888 27436 57916
rect 21416 57876 21422 57888
rect 27430 57876 27436 57888
rect 27488 57916 27494 57928
rect 33410 57916 33416 57928
rect 27488 57888 33416 57916
rect 27488 57876 27494 57888
rect 33410 57876 33416 57888
rect 33468 57876 33474 57928
rect 17862 57808 17868 57860
rect 17920 57848 17926 57860
rect 28442 57848 28448 57860
rect 17920 57820 28448 57848
rect 17920 57808 17926 57820
rect 28442 57808 28448 57820
rect 28500 57808 28506 57860
rect 30558 57848 30564 57860
rect 28966 57820 30564 57848
rect 22830 57740 22836 57792
rect 22888 57780 22894 57792
rect 23934 57780 23940 57792
rect 22888 57752 23940 57780
rect 22888 57740 22894 57752
rect 23934 57740 23940 57752
rect 23992 57740 23998 57792
rect 24762 57740 24768 57792
rect 24820 57780 24826 57792
rect 28966 57780 28994 57820
rect 30558 57808 30564 57820
rect 30616 57808 30622 57860
rect 41414 57808 41420 57860
rect 41472 57848 41478 57860
rect 45922 57848 45928 57860
rect 41472 57820 45928 57848
rect 41472 57808 41478 57820
rect 45922 57808 45928 57820
rect 45980 57808 45986 57860
rect 24820 57752 28994 57780
rect 24820 57740 24826 57752
rect 29178 57740 29184 57792
rect 29236 57780 29242 57792
rect 33962 57780 33968 57792
rect 29236 57752 33968 57780
rect 29236 57740 29242 57752
rect 33962 57740 33968 57752
rect 34020 57740 34026 57792
rect 42886 57740 42892 57792
rect 42944 57780 42950 57792
rect 46842 57780 46848 57792
rect 42944 57752 46848 57780
rect 42944 57740 42950 57752
rect 46842 57740 46848 57752
rect 46900 57780 46906 57792
rect 54110 57780 54116 57792
rect 46900 57752 54116 57780
rect 46900 57740 46906 57752
rect 54110 57740 54116 57752
rect 54168 57740 54174 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 3421 57579 3479 57585
rect 3421 57545 3433 57579
rect 3467 57576 3479 57579
rect 3694 57576 3700 57588
rect 3467 57548 3700 57576
rect 3467 57545 3479 57548
rect 3421 57539 3479 57545
rect 3694 57536 3700 57548
rect 3752 57576 3758 57588
rect 3752 57548 4108 57576
rect 3752 57536 3758 57548
rect 4080 57517 4108 57548
rect 5074 57536 5080 57588
rect 5132 57576 5138 57588
rect 5261 57579 5319 57585
rect 5261 57576 5273 57579
rect 5132 57548 5273 57576
rect 5132 57536 5138 57548
rect 5261 57545 5273 57548
rect 5307 57545 5319 57579
rect 5261 57539 5319 57545
rect 10594 57536 10600 57588
rect 10652 57576 10658 57588
rect 10781 57579 10839 57585
rect 10781 57576 10793 57579
rect 10652 57548 10793 57576
rect 10652 57536 10658 57548
rect 10781 57545 10793 57548
rect 10827 57545 10839 57579
rect 10781 57539 10839 57545
rect 11974 57536 11980 57588
rect 12032 57576 12038 57588
rect 12161 57579 12219 57585
rect 12161 57576 12173 57579
rect 12032 57548 12173 57576
rect 12032 57536 12038 57548
rect 12161 57545 12173 57548
rect 12207 57545 12219 57579
rect 12161 57539 12219 57545
rect 13354 57536 13360 57588
rect 13412 57576 13418 57588
rect 13541 57579 13599 57585
rect 13541 57576 13553 57579
rect 13412 57548 13553 57576
rect 13412 57536 13418 57548
rect 13541 57545 13553 57548
rect 13587 57545 13599 57579
rect 13541 57539 13599 57545
rect 14734 57536 14740 57588
rect 14792 57576 14798 57588
rect 14921 57579 14979 57585
rect 14921 57576 14933 57579
rect 14792 57548 14933 57576
rect 14792 57536 14798 57548
rect 14921 57545 14933 57548
rect 14967 57545 14979 57579
rect 14921 57539 14979 57545
rect 16114 57536 16120 57588
rect 16172 57576 16178 57588
rect 16945 57579 17003 57585
rect 16945 57576 16957 57579
rect 16172 57548 16957 57576
rect 16172 57536 16178 57548
rect 16945 57545 16957 57548
rect 16991 57545 17003 57579
rect 16945 57539 17003 57545
rect 17494 57536 17500 57588
rect 17552 57576 17558 57588
rect 17681 57579 17739 57585
rect 17681 57576 17693 57579
rect 17552 57548 17693 57576
rect 17552 57536 17558 57548
rect 17681 57545 17693 57548
rect 17727 57545 17739 57579
rect 17681 57539 17739 57545
rect 19334 57536 19340 57588
rect 19392 57576 19398 57588
rect 19521 57579 19579 57585
rect 19521 57576 19533 57579
rect 19392 57548 19533 57576
rect 19392 57536 19398 57548
rect 19521 57545 19533 57548
rect 19567 57545 19579 57579
rect 19521 57539 19579 57545
rect 20254 57536 20260 57588
rect 20312 57576 20318 57588
rect 20441 57579 20499 57585
rect 20441 57576 20453 57579
rect 20312 57548 20453 57576
rect 20312 57536 20318 57548
rect 20441 57545 20453 57548
rect 20487 57545 20499 57579
rect 22186 57576 22192 57588
rect 20441 57539 20499 57545
rect 20548 57548 22192 57576
rect 4065 57511 4123 57517
rect 4065 57477 4077 57511
rect 4111 57477 4123 57511
rect 20548 57508 20576 57548
rect 22186 57536 22192 57548
rect 22244 57536 22250 57588
rect 22281 57579 22339 57585
rect 22281 57545 22293 57579
rect 22327 57576 22339 57579
rect 23014 57576 23020 57588
rect 22327 57548 23020 57576
rect 22327 57545 22339 57548
rect 22281 57539 22339 57545
rect 23014 57536 23020 57548
rect 23072 57536 23078 57588
rect 25038 57576 25044 57588
rect 23124 57548 25044 57576
rect 23124 57508 23152 57548
rect 25038 57536 25044 57548
rect 25096 57536 25102 57588
rect 25774 57536 25780 57588
rect 25832 57576 25838 57588
rect 26053 57579 26111 57585
rect 26053 57576 26065 57579
rect 25832 57548 26065 57576
rect 25832 57536 25838 57548
rect 26053 57545 26065 57548
rect 26099 57545 26111 57579
rect 26053 57539 26111 57545
rect 27154 57536 27160 57588
rect 27212 57576 27218 57588
rect 27433 57579 27491 57585
rect 27433 57576 27445 57579
rect 27212 57548 27445 57576
rect 27212 57536 27218 57548
rect 27433 57545 27445 57548
rect 27479 57545 27491 57579
rect 27433 57539 27491 57545
rect 28534 57536 28540 57588
rect 28592 57576 28598 57588
rect 28721 57579 28779 57585
rect 28721 57576 28733 57579
rect 28592 57548 28733 57576
rect 28592 57536 28598 57548
rect 28721 57545 28733 57548
rect 28767 57545 28779 57579
rect 34514 57576 34520 57588
rect 28721 57539 28779 57545
rect 31680 57548 34520 57576
rect 4065 57471 4123 57477
rect 15120 57480 20576 57508
rect 20640 57480 23152 57508
rect 5445 57443 5503 57449
rect 5445 57409 5457 57443
rect 5491 57409 5503 57443
rect 5445 57403 5503 57409
rect 7285 57443 7343 57449
rect 7285 57409 7297 57443
rect 7331 57440 7343 57443
rect 7374 57440 7380 57452
rect 7331 57412 7380 57440
rect 7331 57409 7343 57412
rect 7285 57403 7343 57409
rect 5460 57372 5488 57403
rect 7374 57400 7380 57412
rect 7432 57400 7438 57452
rect 7745 57443 7803 57449
rect 7745 57409 7757 57443
rect 7791 57440 7803 57443
rect 7834 57440 7840 57452
rect 7791 57412 7840 57440
rect 7791 57409 7803 57412
rect 7745 57403 7803 57409
rect 7834 57400 7840 57412
rect 7892 57400 7898 57452
rect 8573 57443 8631 57449
rect 8573 57409 8585 57443
rect 8619 57440 8631 57443
rect 8754 57440 8760 57452
rect 8619 57412 8760 57440
rect 8619 57409 8631 57412
rect 8573 57403 8631 57409
rect 8754 57400 8760 57412
rect 8812 57400 8818 57452
rect 9214 57400 9220 57452
rect 9272 57440 9278 57452
rect 9309 57443 9367 57449
rect 9309 57440 9321 57443
rect 9272 57412 9321 57440
rect 9272 57400 9278 57412
rect 9309 57409 9321 57412
rect 9355 57409 9367 57443
rect 9309 57403 9367 57409
rect 10045 57443 10103 57449
rect 10045 57409 10057 57443
rect 10091 57440 10103 57443
rect 10134 57440 10140 57452
rect 10091 57412 10140 57440
rect 10091 57409 10103 57412
rect 10045 57403 10103 57409
rect 10134 57400 10140 57412
rect 10192 57400 10198 57452
rect 10962 57440 10968 57452
rect 10923 57412 10968 57440
rect 10962 57400 10968 57412
rect 11020 57400 11026 57452
rect 12342 57440 12348 57452
rect 12303 57412 12348 57440
rect 12342 57400 12348 57412
rect 12400 57400 12406 57452
rect 12805 57443 12863 57449
rect 12805 57409 12817 57443
rect 12851 57440 12863 57443
rect 12894 57440 12900 57452
rect 12851 57412 12900 57440
rect 12851 57409 12863 57412
rect 12805 57403 12863 57409
rect 12894 57400 12900 57412
rect 12952 57400 12958 57452
rect 15120 57449 15148 57480
rect 13725 57443 13783 57449
rect 13725 57409 13737 57443
rect 13771 57409 13783 57443
rect 13725 57403 13783 57409
rect 15105 57443 15163 57449
rect 15105 57409 15117 57443
rect 15151 57409 15163 57443
rect 15105 57403 15163 57409
rect 5997 57375 6055 57381
rect 5997 57372 6009 57375
rect 5460 57344 6009 57372
rect 5997 57341 6009 57344
rect 6043 57372 6055 57375
rect 6086 57372 6092 57384
rect 6043 57344 6092 57372
rect 6043 57341 6055 57344
rect 5997 57335 6055 57341
rect 6086 57332 6092 57344
rect 6144 57332 6150 57384
rect 4249 57307 4307 57313
rect 4249 57273 4261 57307
rect 4295 57304 4307 57307
rect 5442 57304 5448 57316
rect 4295 57276 5448 57304
rect 4295 57273 4307 57276
rect 4249 57267 4307 57273
rect 5442 57264 5448 57276
rect 5500 57264 5506 57316
rect 13740 57304 13768 57403
rect 15654 57400 15660 57452
rect 15712 57440 15718 57452
rect 15749 57443 15807 57449
rect 15749 57440 15761 57443
rect 15712 57412 15761 57440
rect 15712 57400 15718 57412
rect 15749 57409 15761 57412
rect 15795 57409 15807 57443
rect 17126 57440 17132 57452
rect 17087 57412 17132 57440
rect 15749 57403 15807 57409
rect 17126 57400 17132 57412
rect 17184 57400 17190 57452
rect 17862 57440 17868 57452
rect 17823 57412 17868 57440
rect 17862 57400 17868 57412
rect 17920 57400 17926 57452
rect 18414 57400 18420 57452
rect 18472 57440 18478 57452
rect 20640 57449 20668 57480
rect 23474 57468 23480 57520
rect 23532 57508 23538 57520
rect 24394 57508 24400 57520
rect 23532 57480 24400 57508
rect 23532 57468 23538 57480
rect 24394 57468 24400 57480
rect 24452 57468 24458 57520
rect 29178 57508 29184 57520
rect 24872 57480 29184 57508
rect 18509 57443 18567 57449
rect 18509 57440 18521 57443
rect 18472 57412 18521 57440
rect 18472 57400 18478 57412
rect 18509 57409 18521 57412
rect 18555 57409 18567 57443
rect 18509 57403 18567 57409
rect 19705 57443 19763 57449
rect 19705 57409 19717 57443
rect 19751 57409 19763 57443
rect 19705 57403 19763 57409
rect 20625 57443 20683 57449
rect 20625 57409 20637 57443
rect 20671 57409 20683 57443
rect 20625 57403 20683 57409
rect 22465 57443 22523 57449
rect 22465 57409 22477 57443
rect 22511 57440 22523 57443
rect 23198 57440 23204 57452
rect 22511 57412 23060 57440
rect 23159 57412 23204 57440
rect 22511 57409 22523 57412
rect 22465 57403 22523 57409
rect 19720 57372 19748 57403
rect 22738 57372 22744 57384
rect 19720 57344 22744 57372
rect 22738 57332 22744 57344
rect 22796 57332 22802 57384
rect 23032 57372 23060 57412
rect 23198 57400 23204 57412
rect 23256 57400 23262 57452
rect 23658 57440 23664 57452
rect 23619 57412 23664 57440
rect 23658 57400 23664 57412
rect 23716 57400 23722 57452
rect 23750 57400 23756 57452
rect 23808 57438 23814 57452
rect 23845 57443 23903 57449
rect 23845 57438 23857 57443
rect 23808 57410 23857 57438
rect 23808 57400 23814 57410
rect 23845 57409 23857 57410
rect 23891 57409 23903 57443
rect 24762 57440 24768 57452
rect 24723 57412 24768 57440
rect 23845 57403 23903 57409
rect 24762 57400 24768 57412
rect 24820 57400 24826 57452
rect 24872 57372 24900 57480
rect 29178 57468 29184 57480
rect 29236 57468 29242 57520
rect 31570 57508 31576 57520
rect 30024 57480 31576 57508
rect 25130 57400 25136 57452
rect 25188 57440 25194 57452
rect 25869 57443 25927 57449
rect 25869 57440 25881 57443
rect 25188 57412 25881 57440
rect 25188 57400 25194 57412
rect 25869 57409 25881 57412
rect 25915 57409 25927 57443
rect 27246 57440 27252 57452
rect 27207 57412 27252 57440
rect 25869 57403 25927 57409
rect 27246 57400 27252 57412
rect 27304 57400 27310 57452
rect 27985 57443 28043 57449
rect 27985 57409 27997 57443
rect 28031 57409 28043 57443
rect 27985 57403 28043 57409
rect 28169 57443 28227 57449
rect 28169 57409 28181 57443
rect 28215 57409 28227 57443
rect 28169 57403 28227 57409
rect 28905 57443 28963 57449
rect 28905 57409 28917 57443
rect 28951 57440 28963 57443
rect 29270 57440 29276 57452
rect 28951 57412 29276 57440
rect 28951 57409 28963 57412
rect 28905 57403 28963 57409
rect 23032 57344 24900 57372
rect 24949 57375 25007 57381
rect 24949 57341 24961 57375
rect 24995 57372 25007 57375
rect 25222 57372 25228 57384
rect 24995 57344 25228 57372
rect 24995 57341 25007 57344
rect 24949 57335 25007 57341
rect 25222 57332 25228 57344
rect 25280 57332 25286 57384
rect 23017 57307 23075 57313
rect 13740 57276 22968 57304
rect 21453 57239 21511 57245
rect 21453 57205 21465 57239
rect 21499 57236 21511 57239
rect 22830 57236 22836 57248
rect 21499 57208 22836 57236
rect 21499 57205 21511 57208
rect 21453 57199 21511 57205
rect 22830 57196 22836 57208
rect 22888 57196 22894 57248
rect 22940 57236 22968 57276
rect 23017 57273 23029 57307
rect 23063 57304 23075 57307
rect 23474 57304 23480 57316
rect 23063 57276 23480 57304
rect 23063 57273 23075 57276
rect 23017 57267 23075 57273
rect 23474 57264 23480 57276
rect 23532 57264 23538 57316
rect 23566 57264 23572 57316
rect 23624 57304 23630 57316
rect 24581 57307 24639 57313
rect 24581 57304 24593 57307
rect 23624 57276 24593 57304
rect 23624 57264 23630 57276
rect 24581 57273 24593 57276
rect 24627 57273 24639 57307
rect 28000 57304 28028 57403
rect 28184 57372 28212 57403
rect 29270 57400 29276 57412
rect 29328 57400 29334 57452
rect 30024 57384 30052 57480
rect 31570 57468 31576 57480
rect 31628 57468 31634 57520
rect 31680 57517 31708 57548
rect 34514 57536 34520 57548
rect 34572 57576 34578 57588
rect 39393 57579 39451 57585
rect 39393 57576 39405 57579
rect 34572 57548 39405 57576
rect 34572 57536 34578 57548
rect 39393 57545 39405 57548
rect 39439 57545 39451 57579
rect 39393 57539 39451 57545
rect 45738 57536 45744 57588
rect 45796 57576 45802 57588
rect 54021 57579 54079 57585
rect 54021 57576 54033 57579
rect 45796 57548 54033 57576
rect 45796 57536 45802 57548
rect 54021 57545 54033 57548
rect 54067 57545 54079 57579
rect 54021 57539 54079 57545
rect 54110 57536 54116 57588
rect 54168 57576 54174 57588
rect 55585 57579 55643 57585
rect 55585 57576 55597 57579
rect 54168 57548 55597 57576
rect 54168 57536 54174 57548
rect 55585 57545 55597 57548
rect 55631 57545 55643 57579
rect 55585 57539 55643 57545
rect 31665 57511 31723 57517
rect 31665 57477 31677 57511
rect 31711 57477 31723 57511
rect 31665 57471 31723 57477
rect 33965 57511 34023 57517
rect 33965 57477 33977 57511
rect 34011 57508 34023 57511
rect 34238 57508 34244 57520
rect 34011 57480 34244 57508
rect 34011 57477 34023 57480
rect 33965 57471 34023 57477
rect 34238 57468 34244 57480
rect 34296 57508 34302 57520
rect 34296 57480 40356 57508
rect 34296 57468 34302 57480
rect 30193 57443 30251 57449
rect 30193 57409 30205 57443
rect 30239 57440 30251 57443
rect 30466 57440 30472 57452
rect 30239 57412 30472 57440
rect 30239 57409 30251 57412
rect 30193 57403 30251 57409
rect 30466 57400 30472 57412
rect 30524 57400 30530 57452
rect 30834 57440 30840 57452
rect 30795 57412 30840 57440
rect 30834 57400 30840 57412
rect 30892 57400 30898 57452
rect 31404 57412 32996 57440
rect 30006 57372 30012 57384
rect 28184 57344 30012 57372
rect 30006 57332 30012 57344
rect 30064 57332 30070 57384
rect 30282 57304 30288 57316
rect 28000 57276 30288 57304
rect 24581 57267 24639 57273
rect 30282 57264 30288 57276
rect 30340 57264 30346 57316
rect 30377 57307 30435 57313
rect 30377 57273 30389 57307
rect 30423 57304 30435 57307
rect 31404 57304 31432 57412
rect 31481 57375 31539 57381
rect 31481 57341 31493 57375
rect 31527 57372 31539 57375
rect 31846 57372 31852 57384
rect 31527 57344 31852 57372
rect 31527 57341 31539 57344
rect 31481 57335 31539 57341
rect 31846 57332 31852 57344
rect 31904 57332 31910 57384
rect 32030 57332 32036 57384
rect 32088 57372 32094 57384
rect 32309 57375 32367 57381
rect 32309 57372 32321 57375
rect 32088 57344 32321 57372
rect 32088 57332 32094 57344
rect 32309 57341 32321 57344
rect 32355 57341 32367 57375
rect 32582 57372 32588 57384
rect 32543 57344 32588 57372
rect 32309 57335 32367 57341
rect 32582 57332 32588 57344
rect 32640 57332 32646 57384
rect 32968 57372 32996 57412
rect 33502 57400 33508 57452
rect 33560 57440 33566 57452
rect 33781 57443 33839 57449
rect 33781 57440 33793 57443
rect 33560 57412 33793 57440
rect 33560 57400 33566 57412
rect 33781 57409 33793 57412
rect 33827 57409 33839 57443
rect 33781 57403 33839 57409
rect 34057 57443 34115 57449
rect 34057 57409 34069 57443
rect 34103 57440 34115 57443
rect 34146 57440 34152 57452
rect 34103 57412 34152 57440
rect 34103 57409 34115 57412
rect 34057 57403 34115 57409
rect 34146 57400 34152 57412
rect 34204 57400 34210 57452
rect 35345 57443 35403 57449
rect 35345 57409 35357 57443
rect 35391 57409 35403 57443
rect 35526 57440 35532 57452
rect 35487 57412 35532 57440
rect 35345 57403 35403 57409
rect 34330 57372 34336 57384
rect 32968 57344 34336 57372
rect 34330 57332 34336 57344
rect 34388 57332 34394 57384
rect 35360 57372 35388 57403
rect 35526 57400 35532 57412
rect 35584 57400 35590 57452
rect 35894 57400 35900 57452
rect 35952 57440 35958 57452
rect 35989 57443 36047 57449
rect 35989 57440 36001 57443
rect 35952 57412 36001 57440
rect 35952 57400 35958 57412
rect 35989 57409 36001 57412
rect 36035 57409 36047 57443
rect 35989 57403 36047 57409
rect 37274 57400 37280 57452
rect 37332 57440 37338 57452
rect 37461 57443 37519 57449
rect 37461 57440 37473 57443
rect 37332 57412 37473 57440
rect 37332 57400 37338 57412
rect 37461 57409 37473 57412
rect 37507 57409 37519 57443
rect 37461 57403 37519 57409
rect 38654 57400 38660 57452
rect 38712 57440 38718 57452
rect 39850 57440 39856 57452
rect 38712 57412 39856 57440
rect 38712 57400 38718 57412
rect 39850 57400 39856 57412
rect 39908 57440 39914 57452
rect 40328 57449 40356 57480
rect 45554 57468 45560 57520
rect 45612 57508 45618 57520
rect 45833 57511 45891 57517
rect 45833 57508 45845 57511
rect 45612 57480 45845 57508
rect 45612 57468 45618 57480
rect 45833 57477 45845 57480
rect 45879 57477 45891 57511
rect 45833 57471 45891 57477
rect 45940 57480 50660 57508
rect 40037 57443 40095 57449
rect 40037 57440 40049 57443
rect 39908 57412 40049 57440
rect 39908 57400 39914 57412
rect 40037 57409 40049 57412
rect 40083 57409 40095 57443
rect 40037 57403 40095 57409
rect 40313 57443 40371 57449
rect 40313 57409 40325 57443
rect 40359 57409 40371 57443
rect 40313 57403 40371 57409
rect 41046 57400 41052 57452
rect 41104 57440 41110 57452
rect 41509 57443 41567 57449
rect 41509 57440 41521 57443
rect 41104 57412 41521 57440
rect 41104 57400 41110 57412
rect 41509 57409 41521 57412
rect 41555 57409 41567 57443
rect 41509 57403 41567 57409
rect 42794 57400 42800 57452
rect 42852 57440 42858 57452
rect 43717 57443 43775 57449
rect 43717 57440 43729 57443
rect 42852 57412 43729 57440
rect 42852 57400 42858 57412
rect 43717 57409 43729 57412
rect 43763 57440 43775 57443
rect 44082 57440 44088 57452
rect 43763 57412 44088 57440
rect 43763 57409 43775 57412
rect 43717 57403 43775 57409
rect 44082 57400 44088 57412
rect 44140 57400 44146 57452
rect 44266 57400 44272 57452
rect 44324 57440 44330 57452
rect 44361 57443 44419 57449
rect 44361 57440 44373 57443
rect 44324 57412 44373 57440
rect 44324 57400 44330 57412
rect 44361 57409 44373 57412
rect 44407 57409 44419 57443
rect 44361 57403 44419 57409
rect 44450 57400 44456 57452
rect 44508 57440 44514 57452
rect 44637 57443 44695 57449
rect 44637 57440 44649 57443
rect 44508 57412 44649 57440
rect 44508 57400 44514 57412
rect 44637 57409 44649 57412
rect 44683 57440 44695 57443
rect 44910 57440 44916 57452
rect 44683 57412 44916 57440
rect 44683 57409 44695 57412
rect 44637 57403 44695 57409
rect 44910 57400 44916 57412
rect 44968 57440 44974 57452
rect 45940 57440 45968 57480
rect 44968 57412 45968 57440
rect 44968 57400 44974 57412
rect 47394 57400 47400 57452
rect 47452 57440 47458 57452
rect 49053 57443 49111 57449
rect 49053 57440 49065 57443
rect 47452 57412 49065 57440
rect 47452 57400 47458 57412
rect 49053 57409 49065 57412
rect 49099 57409 49111 57443
rect 49053 57403 49111 57409
rect 49694 57400 49700 57452
rect 49752 57440 49758 57452
rect 50632 57449 50660 57480
rect 52454 57468 52460 57520
rect 52512 57508 52518 57520
rect 53006 57508 53012 57520
rect 52512 57480 53012 57508
rect 52512 57468 52518 57480
rect 53006 57468 53012 57480
rect 53064 57468 53070 57520
rect 50341 57443 50399 57449
rect 50341 57440 50353 57443
rect 49752 57412 50353 57440
rect 49752 57400 49758 57412
rect 50341 57409 50353 57412
rect 50387 57409 50399 57443
rect 50341 57403 50399 57409
rect 50617 57443 50675 57449
rect 50617 57409 50629 57443
rect 50663 57409 50675 57443
rect 50617 57403 50675 57409
rect 51074 57400 51080 57452
rect 51132 57440 51138 57452
rect 51442 57440 51448 57452
rect 51132 57412 51448 57440
rect 51132 57400 51138 57412
rect 51442 57400 51448 57412
rect 51500 57440 51506 57452
rect 51629 57443 51687 57449
rect 51629 57440 51641 57443
rect 51500 57412 51641 57440
rect 51500 57400 51506 57412
rect 51629 57409 51641 57412
rect 51675 57409 51687 57443
rect 51629 57403 51687 57409
rect 53834 57400 53840 57452
rect 53892 57440 53898 57452
rect 54205 57443 54263 57449
rect 54205 57440 54217 57443
rect 53892 57412 54217 57440
rect 53892 57400 53898 57412
rect 54205 57409 54217 57412
rect 54251 57409 54263 57443
rect 54205 57403 54263 57409
rect 54294 57400 54300 57452
rect 54352 57440 54358 57452
rect 54665 57443 54723 57449
rect 54665 57440 54677 57443
rect 54352 57412 54677 57440
rect 54352 57400 54358 57412
rect 54665 57409 54677 57412
rect 54711 57409 54723 57443
rect 54665 57403 54723 57409
rect 55214 57400 55220 57452
rect 55272 57440 55278 57452
rect 55766 57440 55772 57452
rect 55272 57412 55772 57440
rect 55272 57400 55278 57412
rect 55766 57400 55772 57412
rect 55824 57400 55830 57452
rect 56134 57400 56140 57452
rect 56192 57440 56198 57452
rect 56873 57443 56931 57449
rect 56873 57440 56885 57443
rect 56192 57412 56885 57440
rect 56192 57400 56198 57412
rect 56873 57409 56885 57412
rect 56919 57409 56931 57443
rect 56873 57403 56931 57409
rect 35710 57372 35716 57384
rect 35360 57344 35716 57372
rect 35710 57332 35716 57344
rect 35768 57332 35774 57384
rect 36262 57372 36268 57384
rect 36223 57344 36268 57372
rect 36262 57332 36268 57344
rect 36320 57332 36326 57384
rect 36630 57332 36636 57384
rect 36688 57372 36694 57384
rect 37737 57375 37795 57381
rect 37737 57372 37749 57375
rect 36688 57344 37749 57372
rect 36688 57332 36694 57344
rect 37737 57341 37749 57344
rect 37783 57341 37795 57375
rect 41782 57372 41788 57384
rect 41695 57344 41788 57372
rect 37737 57335 37795 57341
rect 41782 57332 41788 57344
rect 41840 57372 41846 57384
rect 42978 57372 42984 57384
rect 41840 57344 42984 57372
rect 41840 57332 41846 57344
rect 42978 57332 42984 57344
rect 43036 57332 43042 57384
rect 43441 57375 43499 57381
rect 43441 57341 43453 57375
rect 43487 57372 43499 57375
rect 43622 57372 43628 57384
rect 43487 57344 43628 57372
rect 43487 57341 43499 57344
rect 43441 57335 43499 57341
rect 43622 57332 43628 57344
rect 43680 57332 43686 57384
rect 43990 57332 43996 57384
rect 44048 57372 44054 57384
rect 44545 57375 44603 57381
rect 44545 57372 44557 57375
rect 44048 57344 44557 57372
rect 44048 57332 44054 57344
rect 44545 57341 44557 57344
rect 44591 57372 44603 57375
rect 45738 57372 45744 57384
rect 44591 57344 45744 57372
rect 44591 57341 44603 57344
rect 44545 57335 44603 57341
rect 45738 57332 45744 57344
rect 45796 57332 45802 57384
rect 46934 57332 46940 57384
rect 46992 57372 46998 57384
rect 47765 57375 47823 57381
rect 47765 57372 47777 57375
rect 46992 57344 47777 57372
rect 46992 57332 46998 57344
rect 47765 57341 47777 57344
rect 47811 57341 47823 57375
rect 47765 57335 47823 57341
rect 35161 57307 35219 57313
rect 35161 57304 35173 57307
rect 30423 57276 31432 57304
rect 31496 57276 35173 57304
rect 30423 57273 30435 57276
rect 30377 57267 30435 57273
rect 23842 57236 23848 57248
rect 22940 57208 23848 57236
rect 23842 57196 23848 57208
rect 23900 57196 23906 57248
rect 24026 57236 24032 57248
rect 23987 57208 24032 57236
rect 24026 57196 24032 57208
rect 24084 57196 24090 57248
rect 24118 57196 24124 57248
rect 24176 57236 24182 57248
rect 25314 57236 25320 57248
rect 24176 57208 25320 57236
rect 24176 57196 24182 57208
rect 25314 57196 25320 57208
rect 25372 57196 25378 57248
rect 28169 57239 28227 57245
rect 28169 57205 28181 57239
rect 28215 57236 28227 57239
rect 28810 57236 28816 57248
rect 28215 57208 28816 57236
rect 28215 57205 28227 57208
rect 28169 57199 28227 57205
rect 28810 57196 28816 57208
rect 28868 57196 28874 57248
rect 28902 57196 28908 57248
rect 28960 57236 28966 57248
rect 31496 57236 31524 57276
rect 35161 57273 35173 57276
rect 35207 57273 35219 57307
rect 35161 57267 35219 57273
rect 36722 57264 36728 57316
rect 36780 57304 36786 57316
rect 38930 57304 38936 57316
rect 36780 57276 38936 57304
rect 36780 57264 36786 57276
rect 38930 57264 38936 57276
rect 38988 57304 38994 57316
rect 40678 57304 40684 57316
rect 38988 57276 40684 57304
rect 38988 57264 38994 57276
rect 40678 57264 40684 57276
rect 40736 57264 40742 57316
rect 41230 57264 41236 57316
rect 41288 57304 41294 57316
rect 41693 57307 41751 57313
rect 41693 57304 41705 57307
rect 41288 57276 41705 57304
rect 41288 57264 41294 57276
rect 41693 57273 41705 57276
rect 41739 57273 41751 57307
rect 41693 57267 41751 57273
rect 45646 57264 45652 57316
rect 45704 57304 45710 57316
rect 47780 57304 47808 57335
rect 55674 57332 55680 57384
rect 55732 57372 55738 57384
rect 56229 57375 56287 57381
rect 56229 57372 56241 57375
rect 55732 57344 56241 57372
rect 55732 57332 55738 57344
rect 56229 57341 56241 57344
rect 56275 57341 56287 57375
rect 56229 57335 56287 57341
rect 49697 57307 49755 57313
rect 49697 57304 49709 57307
rect 45704 57276 47164 57304
rect 47780 57276 49709 57304
rect 45704 57264 45710 57276
rect 28960 57208 31524 57236
rect 28960 57196 28966 57208
rect 31570 57196 31576 57248
rect 31628 57236 31634 57248
rect 33597 57239 33655 57245
rect 33597 57236 33609 57239
rect 31628 57208 33609 57236
rect 31628 57196 31634 57208
rect 33597 57205 33609 57208
rect 33643 57205 33655 57239
rect 38746 57236 38752 57248
rect 38707 57208 38752 57236
rect 33597 57199 33655 57205
rect 38746 57196 38752 57208
rect 38804 57196 38810 57248
rect 40494 57196 40500 57248
rect 40552 57236 40558 57248
rect 41325 57239 41383 57245
rect 41325 57236 41337 57239
rect 40552 57208 41337 57236
rect 40552 57196 40558 57208
rect 41325 57205 41337 57208
rect 41371 57205 41383 57239
rect 41325 57199 41383 57205
rect 43346 57196 43352 57248
rect 43404 57236 43410 57248
rect 44177 57239 44235 57245
rect 44177 57236 44189 57239
rect 43404 57208 44189 57236
rect 43404 57196 43410 57208
rect 44177 57205 44189 57208
rect 44223 57205 44235 57239
rect 44177 57199 44235 57205
rect 45462 57196 45468 57248
rect 45520 57236 45526 57248
rect 45741 57239 45799 57245
rect 45741 57236 45753 57239
rect 45520 57208 45753 57236
rect 45520 57196 45526 57208
rect 45741 57205 45753 57208
rect 45787 57205 45799 57239
rect 46382 57236 46388 57248
rect 46343 57208 46388 57236
rect 45741 57199 45799 57205
rect 46382 57196 46388 57208
rect 46440 57196 46446 57248
rect 47026 57236 47032 57248
rect 46987 57208 47032 57236
rect 47026 57196 47032 57208
rect 47084 57196 47090 57248
rect 47136 57236 47164 57276
rect 49697 57273 49709 57276
rect 49743 57273 49755 57307
rect 49697 57267 49755 57273
rect 47995 57239 48053 57245
rect 47995 57236 48007 57239
rect 47136 57208 48007 57236
rect 47995 57205 48007 57208
rect 48041 57205 48053 57239
rect 51810 57236 51816 57248
rect 51771 57208 51816 57236
rect 47995 57199 48053 57205
rect 51810 57196 51816 57208
rect 51868 57196 51874 57248
rect 53098 57236 53104 57248
rect 53059 57208 53104 57236
rect 53098 57196 53104 57208
rect 53156 57196 53162 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 4614 56992 4620 57044
rect 4672 57032 4678 57044
rect 4709 57035 4767 57041
rect 4709 57032 4721 57035
rect 4672 57004 4721 57032
rect 4672 56992 4678 57004
rect 4709 57001 4721 57004
rect 4755 57001 4767 57035
rect 4709 56995 4767 57001
rect 5905 57035 5963 57041
rect 5905 57001 5917 57035
rect 5951 57032 5963 57035
rect 5994 57032 6000 57044
rect 5951 57004 6000 57032
rect 5951 57001 5963 57004
rect 5905 56995 5963 57001
rect 5994 56992 6000 57004
rect 6052 56992 6058 57044
rect 6454 56992 6460 57044
rect 6512 57032 6518 57044
rect 6549 57035 6607 57041
rect 6549 57032 6561 57035
rect 6512 57004 6561 57032
rect 6512 56992 6518 57004
rect 6549 57001 6561 57004
rect 6595 57001 6607 57035
rect 6549 56995 6607 57001
rect 11514 56992 11520 57044
rect 11572 57032 11578 57044
rect 11609 57035 11667 57041
rect 11609 57032 11621 57035
rect 11572 57004 11621 57032
rect 11572 56992 11578 57004
rect 11609 57001 11621 57004
rect 11655 57001 11667 57035
rect 11609 56995 11667 57001
rect 14274 56992 14280 57044
rect 14332 57032 14338 57044
rect 14369 57035 14427 57041
rect 14369 57032 14381 57035
rect 14332 57004 14381 57032
rect 14332 56992 14338 57004
rect 14369 57001 14381 57004
rect 14415 57001 14427 57035
rect 14369 56995 14427 57001
rect 17034 56992 17040 57044
rect 17092 57032 17098 57044
rect 17129 57035 17187 57041
rect 17129 57032 17141 57035
rect 17092 57004 17141 57032
rect 17092 56992 17098 57004
rect 17129 57001 17141 57004
rect 17175 57001 17187 57035
rect 17129 56995 17187 57001
rect 19889 57035 19947 57041
rect 19889 57001 19901 57035
rect 19935 57032 19947 57035
rect 19978 57032 19984 57044
rect 19935 57004 19984 57032
rect 19935 57001 19947 57004
rect 19889 56995 19947 57001
rect 19978 56992 19984 57004
rect 20036 56992 20042 57044
rect 21085 57035 21143 57041
rect 21085 57001 21097 57035
rect 21131 57032 21143 57035
rect 21174 57032 21180 57044
rect 21131 57004 21180 57032
rect 21131 57001 21143 57004
rect 21085 56995 21143 57001
rect 21174 56992 21180 57004
rect 21232 56992 21238 57044
rect 21634 56992 21640 57044
rect 21692 57032 21698 57044
rect 21821 57035 21879 57041
rect 21821 57032 21833 57035
rect 21692 57004 21833 57032
rect 21692 56992 21698 57004
rect 21821 57001 21833 57004
rect 21867 57001 21879 57035
rect 21821 56995 21879 57001
rect 23198 56992 23204 57044
rect 23256 57032 23262 57044
rect 23477 57035 23535 57041
rect 23477 57032 23489 57035
rect 23256 57004 23489 57032
rect 23256 56992 23262 57004
rect 23477 57001 23489 57004
rect 23523 57001 23535 57035
rect 23477 56995 23535 57001
rect 23842 56992 23848 57044
rect 23900 57032 23906 57044
rect 24029 57035 24087 57041
rect 24029 57032 24041 57035
rect 23900 57004 24041 57032
rect 23900 56992 23906 57004
rect 24029 57001 24041 57004
rect 24075 57001 24087 57035
rect 24029 56995 24087 57001
rect 27154 56992 27160 57044
rect 27212 57032 27218 57044
rect 27249 57035 27307 57041
rect 27249 57032 27261 57035
rect 27212 57004 27261 57032
rect 27212 56992 27218 57004
rect 27249 57001 27261 57004
rect 27295 57001 27307 57035
rect 27249 56995 27307 57001
rect 27430 56992 27436 57044
rect 27488 57032 27494 57044
rect 27614 57032 27620 57044
rect 27488 57004 27620 57032
rect 27488 56992 27494 57004
rect 27614 56992 27620 57004
rect 27672 56992 27678 57044
rect 27709 57035 27767 57041
rect 27709 57001 27721 57035
rect 27755 57032 27767 57035
rect 28902 57032 28908 57044
rect 27755 57004 28908 57032
rect 27755 57001 27767 57004
rect 27709 56995 27767 57001
rect 28902 56992 28908 57004
rect 28960 56992 28966 57044
rect 31294 57032 31300 57044
rect 31255 57004 31300 57032
rect 31294 56992 31300 57004
rect 31352 56992 31358 57044
rect 36446 57032 36452 57044
rect 31404 57004 36452 57032
rect 10962 56924 10968 56976
rect 11020 56964 11026 56976
rect 11149 56967 11207 56973
rect 11149 56964 11161 56967
rect 11020 56936 11161 56964
rect 11020 56924 11026 56936
rect 11149 56933 11161 56936
rect 11195 56964 11207 56967
rect 21358 56964 21364 56976
rect 11195 56936 21364 56964
rect 11195 56933 11207 56936
rect 11149 56927 11207 56933
rect 21358 56924 21364 56936
rect 21416 56924 21422 56976
rect 22925 56967 22983 56973
rect 22925 56933 22937 56967
rect 22971 56964 22983 56967
rect 24118 56964 24124 56976
rect 22971 56936 24124 56964
rect 22971 56933 22983 56936
rect 22925 56927 22983 56933
rect 24118 56924 24124 56936
rect 24176 56924 24182 56976
rect 28350 56964 28356 56976
rect 26620 56936 28356 56964
rect 22738 56856 22744 56908
rect 22796 56896 22802 56908
rect 23385 56899 23443 56905
rect 23385 56896 23397 56899
rect 22796 56868 23397 56896
rect 22796 56856 22802 56868
rect 23385 56865 23397 56868
rect 23431 56896 23443 56899
rect 23750 56896 23756 56908
rect 23431 56868 23756 56896
rect 23431 56865 23443 56868
rect 23385 56859 23443 56865
rect 23750 56856 23756 56868
rect 23808 56856 23814 56908
rect 25038 56896 25044 56908
rect 24999 56868 25044 56896
rect 25038 56856 25044 56868
rect 25096 56856 25102 56908
rect 22005 56831 22063 56837
rect 22005 56797 22017 56831
rect 22051 56828 22063 56831
rect 23474 56828 23480 56840
rect 22051 56800 23480 56828
rect 22051 56797 22063 56800
rect 22005 56791 22063 56797
rect 23474 56788 23480 56800
rect 23532 56788 23538 56840
rect 23891 56831 23949 56837
rect 23891 56797 23903 56831
rect 23937 56828 23949 56831
rect 24762 56828 24768 56840
rect 23937 56800 24768 56828
rect 23937 56797 23949 56800
rect 23891 56791 23949 56797
rect 24762 56788 24768 56800
rect 24820 56788 24826 56840
rect 25130 56788 25136 56840
rect 25188 56828 25194 56840
rect 25504 56831 25562 56837
rect 25188 56800 25233 56828
rect 25188 56788 25194 56800
rect 25504 56797 25516 56831
rect 25550 56828 25562 56831
rect 25682 56828 25688 56840
rect 25550 56800 25688 56828
rect 25550 56797 25562 56800
rect 25504 56791 25562 56797
rect 25682 56788 25688 56800
rect 25740 56788 25746 56840
rect 26620 56837 26648 56936
rect 28350 56924 28356 56936
rect 28408 56924 28414 56976
rect 28442 56924 28448 56976
rect 28500 56964 28506 56976
rect 28537 56967 28595 56973
rect 28537 56964 28549 56967
rect 28500 56936 28549 56964
rect 28500 56924 28506 56936
rect 28537 56933 28549 56936
rect 28583 56933 28595 56967
rect 28810 56964 28816 56976
rect 28771 56936 28816 56964
rect 28537 56927 28595 56933
rect 28810 56924 28816 56936
rect 28868 56924 28874 56976
rect 31404 56964 31432 57004
rect 36446 56992 36452 57004
rect 36504 56992 36510 57044
rect 36538 56992 36544 57044
rect 36596 57032 36602 57044
rect 41046 57032 41052 57044
rect 36596 57004 40448 57032
rect 41007 57004 41052 57032
rect 36596 56992 36602 57004
rect 28920 56936 31432 56964
rect 31757 56967 31815 56973
rect 28258 56896 28264 56908
rect 26804 56868 28264 56896
rect 26804 56837 26832 56868
rect 28258 56856 28264 56868
rect 28316 56896 28322 56908
rect 28316 56868 28856 56896
rect 28316 56856 28322 56868
rect 26605 56831 26663 56837
rect 26605 56797 26617 56831
rect 26651 56797 26663 56831
rect 26605 56791 26663 56797
rect 26789 56831 26847 56837
rect 26789 56797 26801 56831
rect 26835 56797 26847 56831
rect 27430 56828 27436 56840
rect 27391 56800 27436 56828
rect 26789 56791 26847 56797
rect 27430 56788 27436 56800
rect 27488 56788 27494 56840
rect 27522 56788 27528 56840
rect 27580 56828 27586 56840
rect 27798 56828 27804 56840
rect 27580 56800 27625 56828
rect 27759 56800 27804 56828
rect 27580 56788 27586 56800
rect 27798 56788 27804 56800
rect 27856 56788 27862 56840
rect 28721 56831 28779 56837
rect 28721 56797 28733 56831
rect 28767 56797 28779 56831
rect 28721 56791 28779 56797
rect 22186 56720 22192 56772
rect 22244 56760 22250 56772
rect 26697 56763 26755 56769
rect 22244 56732 25728 56760
rect 22244 56720 22250 56732
rect 23842 56692 23848 56704
rect 23803 56664 23848 56692
rect 23842 56652 23848 56664
rect 23900 56652 23906 56704
rect 25501 56695 25559 56701
rect 25501 56661 25513 56695
rect 25547 56692 25559 56695
rect 25590 56692 25596 56704
rect 25547 56664 25596 56692
rect 25547 56661 25559 56664
rect 25501 56655 25559 56661
rect 25590 56652 25596 56664
rect 25648 56652 25654 56704
rect 25700 56701 25728 56732
rect 26697 56729 26709 56763
rect 26743 56760 26755 56763
rect 28736 56760 28764 56791
rect 26743 56732 28764 56760
rect 26743 56729 26755 56732
rect 26697 56723 26755 56729
rect 25685 56695 25743 56701
rect 25685 56661 25697 56695
rect 25731 56661 25743 56695
rect 25685 56655 25743 56661
rect 27522 56652 27528 56704
rect 27580 56692 27586 56704
rect 28718 56692 28724 56704
rect 27580 56664 28724 56692
rect 27580 56652 27586 56664
rect 28718 56652 28724 56664
rect 28776 56652 28782 56704
rect 28828 56692 28856 56868
rect 28920 56837 28948 56936
rect 31757 56933 31769 56967
rect 31803 56933 31815 56967
rect 31757 56927 31815 56933
rect 28997 56899 29055 56905
rect 28997 56865 29009 56899
rect 29043 56896 29055 56899
rect 29270 56896 29276 56908
rect 29043 56868 29276 56896
rect 29043 56865 29055 56868
rect 28997 56859 29055 56865
rect 29270 56856 29276 56868
rect 29328 56896 29334 56908
rect 29733 56899 29791 56905
rect 29733 56896 29745 56899
rect 29328 56868 29745 56896
rect 29328 56856 29334 56868
rect 29733 56865 29745 56868
rect 29779 56865 29791 56899
rect 29733 56859 29791 56865
rect 30006 56856 30012 56908
rect 30064 56896 30070 56908
rect 30193 56899 30251 56905
rect 30193 56896 30205 56899
rect 30064 56868 30205 56896
rect 30064 56856 30070 56868
rect 30193 56865 30205 56868
rect 30239 56865 30251 56899
rect 31772 56896 31800 56927
rect 31938 56924 31944 56976
rect 31996 56964 32002 56976
rect 33229 56967 33287 56973
rect 33229 56964 33241 56967
rect 31996 56936 33241 56964
rect 31996 56924 32002 56936
rect 33229 56933 33241 56936
rect 33275 56933 33287 56967
rect 33229 56927 33287 56933
rect 33962 56924 33968 56976
rect 34020 56964 34026 56976
rect 36357 56967 36415 56973
rect 36357 56964 36369 56967
rect 34020 56936 36369 56964
rect 34020 56924 34026 56936
rect 36357 56933 36369 56936
rect 36403 56933 36415 56967
rect 39301 56967 39359 56973
rect 39301 56964 39313 56967
rect 36357 56927 36415 56933
rect 38120 56936 39313 56964
rect 31772 56868 33088 56896
rect 30193 56859 30251 56865
rect 28905 56831 28963 56837
rect 28905 56797 28917 56831
rect 28951 56797 28963 56831
rect 29178 56828 29184 56840
rect 29139 56800 29184 56828
rect 28905 56791 28963 56797
rect 29178 56788 29184 56800
rect 29236 56788 29242 56840
rect 29917 56831 29975 56837
rect 29917 56797 29929 56831
rect 29963 56828 29975 56831
rect 30101 56831 30159 56837
rect 29963 56800 30052 56828
rect 29963 56797 29975 56800
rect 29917 56791 29975 56797
rect 30024 56772 30052 56800
rect 30101 56797 30113 56831
rect 30147 56797 30159 56831
rect 30282 56828 30288 56840
rect 30243 56800 30288 56828
rect 30101 56791 30159 56797
rect 30006 56720 30012 56772
rect 30064 56720 30070 56772
rect 30116 56692 30144 56791
rect 30282 56788 30288 56800
rect 30340 56788 30346 56840
rect 30374 56788 30380 56840
rect 30432 56828 30438 56840
rect 30469 56831 30527 56837
rect 30469 56828 30481 56831
rect 30432 56800 30481 56828
rect 30432 56788 30438 56800
rect 30469 56797 30481 56800
rect 30515 56797 30527 56831
rect 30469 56791 30527 56797
rect 31846 56788 31852 56840
rect 31904 56837 31910 56840
rect 31904 56831 31940 56837
rect 31928 56797 31940 56831
rect 32306 56828 32312 56840
rect 32267 56800 32312 56828
rect 31904 56791 31940 56797
rect 31904 56788 31910 56791
rect 32306 56788 32312 56800
rect 32364 56788 32370 56840
rect 32401 56831 32459 56837
rect 32401 56797 32413 56831
rect 32447 56828 32459 56831
rect 32950 56828 32956 56840
rect 32447 56800 32956 56828
rect 32447 56797 32459 56800
rect 32401 56791 32459 56797
rect 32950 56788 32956 56800
rect 33008 56788 33014 56840
rect 33060 56837 33088 56868
rect 33410 56856 33416 56908
rect 33468 56896 33474 56908
rect 35069 56899 35127 56905
rect 35069 56896 35081 56899
rect 33468 56868 35081 56896
rect 33468 56856 33474 56868
rect 35069 56865 35081 56868
rect 35115 56865 35127 56899
rect 35069 56859 35127 56865
rect 35253 56899 35311 56905
rect 35253 56865 35265 56899
rect 35299 56896 35311 56899
rect 35526 56896 35532 56908
rect 35299 56868 35532 56896
rect 35299 56865 35311 56868
rect 35253 56859 35311 56865
rect 35526 56856 35532 56868
rect 35584 56896 35590 56908
rect 38013 56899 38071 56905
rect 38013 56896 38025 56899
rect 35584 56868 38025 56896
rect 35584 56856 35590 56868
rect 38013 56865 38025 56868
rect 38059 56865 38071 56899
rect 38013 56859 38071 56865
rect 33045 56831 33103 56837
rect 33045 56797 33057 56831
rect 33091 56797 33103 56831
rect 33045 56791 33103 56797
rect 33226 56788 33232 56840
rect 33284 56828 33290 56840
rect 33321 56831 33379 56837
rect 33321 56828 33333 56831
rect 33284 56800 33333 56828
rect 33284 56788 33290 56800
rect 33321 56797 33333 56800
rect 33367 56797 33379 56831
rect 33962 56828 33968 56840
rect 33923 56800 33968 56828
rect 33321 56791 33379 56797
rect 33962 56788 33968 56800
rect 34020 56788 34026 56840
rect 34146 56828 34152 56840
rect 34059 56800 34152 56828
rect 34146 56788 34152 56800
rect 34204 56788 34210 56840
rect 34238 56788 34244 56840
rect 34296 56828 34302 56840
rect 35437 56831 35495 56837
rect 34296 56800 34341 56828
rect 34296 56788 34302 56800
rect 35437 56797 35449 56831
rect 35483 56797 35495 56831
rect 35437 56791 35495 56797
rect 35621 56831 35679 56837
rect 35621 56797 35633 56831
rect 35667 56828 35679 56831
rect 35986 56828 35992 56840
rect 35667 56800 35992 56828
rect 35667 56797 35679 56800
rect 35621 56791 35679 56797
rect 33781 56763 33839 56769
rect 33781 56760 33793 56763
rect 31726 56732 33793 56760
rect 28828 56664 30144 56692
rect 30282 56652 30288 56704
rect 30340 56692 30346 56704
rect 31726 56692 31754 56732
rect 33781 56729 33793 56732
rect 33827 56729 33839 56763
rect 34164 56760 34192 56788
rect 34882 56760 34888 56772
rect 34164 56732 34888 56760
rect 33781 56723 33839 56729
rect 34882 56720 34888 56732
rect 34940 56720 34946 56772
rect 35452 56760 35480 56791
rect 35986 56788 35992 56800
rect 36044 56828 36050 56840
rect 36265 56831 36323 56837
rect 36265 56828 36277 56831
rect 36044 56800 36277 56828
rect 36044 56788 36050 56800
rect 36265 56797 36277 56800
rect 36311 56797 36323 56831
rect 36538 56828 36544 56840
rect 36499 56800 36544 56828
rect 36265 56791 36323 56797
rect 36538 56788 36544 56800
rect 36596 56788 36602 56840
rect 36722 56828 36728 56840
rect 36683 56800 36728 56828
rect 36722 56788 36728 56800
rect 36780 56788 36786 56840
rect 36906 56788 36912 56840
rect 36964 56828 36970 56840
rect 37001 56831 37059 56837
rect 37001 56828 37013 56831
rect 36964 56800 37013 56828
rect 36964 56788 36970 56800
rect 37001 56797 37013 56800
rect 37047 56797 37059 56831
rect 37001 56791 37059 56797
rect 35710 56760 35716 56772
rect 35452 56732 35716 56760
rect 35710 56720 35716 56732
rect 35768 56760 35774 56772
rect 38120 56760 38148 56936
rect 39301 56933 39313 56936
rect 39347 56933 39359 56967
rect 40420 56964 40448 57004
rect 41046 56992 41052 57004
rect 41104 56992 41110 57044
rect 41601 57035 41659 57041
rect 41601 57001 41613 57035
rect 41647 57032 41659 57035
rect 42702 57032 42708 57044
rect 41647 57004 42708 57032
rect 41647 57001 41659 57004
rect 41601 56995 41659 57001
rect 42702 56992 42708 57004
rect 42760 56992 42766 57044
rect 42886 57032 42892 57044
rect 42847 57004 42892 57032
rect 42886 56992 42892 57004
rect 42944 56992 42950 57044
rect 43254 56992 43260 57044
rect 43312 57032 43318 57044
rect 43312 57004 44864 57032
rect 43312 56992 43318 57004
rect 43441 56967 43499 56973
rect 43441 56964 43453 56967
rect 40420 56936 43453 56964
rect 39301 56927 39359 56933
rect 43441 56933 43453 56936
rect 43487 56933 43499 56967
rect 43441 56927 43499 56933
rect 38197 56899 38255 56905
rect 38197 56865 38209 56899
rect 38243 56896 38255 56899
rect 38654 56896 38660 56908
rect 38243 56868 38660 56896
rect 38243 56865 38255 56868
rect 38197 56859 38255 56865
rect 38654 56856 38660 56868
rect 38712 56896 38718 56908
rect 38712 56868 38884 56896
rect 38712 56856 38718 56868
rect 38289 56831 38347 56837
rect 38289 56797 38301 56831
rect 38335 56797 38347 56831
rect 38289 56791 38347 56797
rect 38381 56831 38439 56837
rect 38381 56797 38393 56831
rect 38427 56797 38439 56831
rect 38381 56791 38439 56797
rect 35768 56732 38148 56760
rect 35768 56720 35774 56732
rect 31938 56692 31944 56704
rect 30340 56664 31754 56692
rect 31899 56664 31944 56692
rect 30340 56652 30346 56664
rect 31938 56652 31944 56664
rect 31996 56652 32002 56704
rect 32306 56652 32312 56704
rect 32364 56692 32370 56704
rect 32861 56695 32919 56701
rect 32861 56692 32873 56695
rect 32364 56664 32873 56692
rect 32364 56652 32370 56664
rect 32861 56661 32873 56664
rect 32907 56661 32919 56695
rect 32861 56655 32919 56661
rect 32950 56652 32956 56704
rect 33008 56692 33014 56704
rect 33502 56692 33508 56704
rect 33008 56664 33508 56692
rect 33008 56652 33014 56664
rect 33502 56652 33508 56664
rect 33560 56652 33566 56704
rect 38304 56692 38332 56791
rect 38396 56760 38424 56791
rect 38470 56788 38476 56840
rect 38528 56828 38534 56840
rect 38856 56828 38884 56868
rect 40126 56856 40132 56908
rect 40184 56896 40190 56908
rect 40313 56899 40371 56905
rect 40313 56896 40325 56899
rect 40184 56868 40325 56896
rect 40184 56856 40190 56868
rect 40313 56865 40325 56868
rect 40359 56865 40371 56899
rect 40494 56896 40500 56908
rect 40455 56868 40500 56896
rect 40313 56859 40371 56865
rect 40494 56856 40500 56868
rect 40552 56856 40558 56908
rect 40678 56856 40684 56908
rect 40736 56896 40742 56908
rect 41693 56899 41751 56905
rect 41693 56896 41705 56899
rect 40736 56868 41705 56896
rect 40736 56856 40742 56868
rect 41693 56865 41705 56868
rect 41739 56896 41751 56899
rect 43346 56896 43352 56908
rect 41739 56868 42472 56896
rect 43307 56868 43352 56896
rect 41739 56865 41751 56868
rect 41693 56859 41751 56865
rect 39025 56831 39083 56837
rect 39025 56828 39037 56831
rect 38528 56800 38573 56828
rect 38856 56800 39037 56828
rect 38528 56788 38534 56800
rect 39025 56797 39037 56800
rect 39071 56797 39083 56831
rect 39025 56791 39083 56797
rect 40218 56788 40224 56840
rect 40276 56828 40282 56840
rect 40405 56831 40463 56837
rect 40276 56800 40321 56828
rect 40276 56788 40282 56800
rect 40405 56797 40417 56831
rect 40451 56828 40463 56831
rect 41174 56831 41232 56837
rect 41174 56828 41186 56831
rect 40451 56800 41186 56828
rect 40451 56797 40463 56800
rect 40405 56791 40463 56797
rect 41174 56797 41186 56800
rect 41220 56828 41232 56831
rect 41782 56828 41788 56840
rect 41220 56800 41788 56828
rect 41220 56797 41232 56800
rect 41174 56791 41232 56797
rect 41782 56788 41788 56800
rect 41840 56788 41846 56840
rect 42150 56828 42156 56840
rect 42111 56800 42156 56828
rect 42150 56788 42156 56800
rect 42208 56788 42214 56840
rect 42444 56828 42472 56868
rect 43346 56856 43352 56868
rect 43404 56856 43410 56908
rect 44358 56896 44364 56908
rect 43916 56868 44364 56896
rect 43070 56828 43076 56840
rect 42444 56800 43076 56828
rect 43070 56788 43076 56800
rect 43128 56828 43134 56840
rect 43916 56837 43944 56868
rect 44358 56856 44364 56868
rect 44416 56856 44422 56908
rect 44836 56896 44864 57004
rect 46014 56992 46020 57044
rect 46072 57032 46078 57044
rect 47765 57035 47823 57041
rect 47765 57032 47777 57035
rect 46072 57004 47777 57032
rect 46072 56992 46078 57004
rect 47765 57001 47777 57004
rect 47811 57001 47823 57035
rect 47765 56995 47823 57001
rect 50154 56992 50160 57044
rect 50212 57032 50218 57044
rect 50341 57035 50399 57041
rect 50341 57032 50353 57035
rect 50212 57004 50353 57032
rect 50212 56992 50218 57004
rect 50341 57001 50353 57004
rect 50387 57001 50399 57035
rect 50341 56995 50399 57001
rect 50614 56992 50620 57044
rect 50672 57032 50678 57044
rect 50985 57035 51043 57041
rect 50985 57032 50997 57035
rect 50672 57004 50997 57032
rect 50672 56992 50678 57004
rect 50985 57001 50997 57004
rect 51031 57001 51043 57035
rect 50985 56995 51043 57001
rect 51534 56992 51540 57044
rect 51592 57032 51598 57044
rect 51629 57035 51687 57041
rect 51629 57032 51641 57035
rect 51592 57004 51641 57032
rect 51592 56992 51598 57004
rect 51629 57001 51641 57004
rect 51675 57001 51687 57035
rect 51629 56995 51687 57001
rect 51994 56992 52000 57044
rect 52052 57032 52058 57044
rect 52273 57035 52331 57041
rect 52273 57032 52285 57035
rect 52052 57004 52285 57032
rect 52052 56992 52058 57004
rect 52273 57001 52285 57004
rect 52319 57001 52331 57035
rect 52273 56995 52331 57001
rect 52914 56992 52920 57044
rect 52972 57032 52978 57044
rect 53009 57035 53067 57041
rect 53009 57032 53021 57035
rect 52972 57004 53021 57032
rect 52972 56992 52978 57004
rect 53009 57001 53021 57004
rect 53055 57001 53067 57035
rect 53009 56995 53067 57001
rect 53374 56992 53380 57044
rect 53432 57032 53438 57044
rect 53653 57035 53711 57041
rect 53653 57032 53665 57035
rect 53432 57004 53665 57032
rect 53432 56992 53438 57004
rect 53653 57001 53665 57004
rect 53699 57001 53711 57035
rect 53653 56995 53711 57001
rect 53834 56992 53840 57044
rect 53892 57032 53898 57044
rect 54297 57035 54355 57041
rect 54297 57032 54309 57035
rect 53892 57004 54309 57032
rect 53892 56992 53898 57004
rect 54297 57001 54309 57004
rect 54343 57001 54355 57035
rect 54297 56995 54355 57001
rect 55766 56992 55772 57044
rect 55824 57032 55830 57044
rect 56137 57035 56195 57041
rect 56137 57032 56149 57035
rect 55824 57004 56149 57032
rect 55824 56992 55830 57004
rect 56137 57001 56149 57004
rect 56183 57001 56195 57035
rect 56137 56995 56195 57001
rect 45094 56924 45100 56976
rect 45152 56964 45158 56976
rect 47121 56967 47179 56973
rect 47121 56964 47133 56967
rect 45152 56936 47133 56964
rect 45152 56924 45158 56936
rect 47121 56933 47133 56936
rect 47167 56933 47179 56967
rect 47121 56927 47179 56933
rect 46477 56899 46535 56905
rect 46477 56896 46489 56899
rect 44836 56868 46489 56896
rect 46477 56865 46489 56868
rect 46523 56865 46535 56899
rect 46477 56859 46535 56865
rect 48314 56856 48320 56908
rect 48372 56896 48378 56908
rect 48409 56899 48467 56905
rect 48409 56896 48421 56899
rect 48372 56868 48421 56896
rect 48372 56856 48378 56868
rect 48409 56865 48421 56868
rect 48455 56896 48467 56899
rect 49697 56899 49755 56905
rect 49697 56896 49709 56899
rect 48455 56868 49709 56896
rect 48455 56865 48467 56868
rect 48409 56859 48467 56865
rect 49697 56865 49709 56868
rect 49743 56865 49755 56899
rect 49697 56859 49755 56865
rect 43533 56831 43591 56837
rect 43533 56828 43545 56831
rect 43128 56800 43545 56828
rect 43128 56788 43134 56800
rect 43533 56797 43545 56800
rect 43579 56797 43591 56831
rect 43533 56791 43591 56797
rect 43901 56831 43959 56837
rect 43901 56797 43913 56831
rect 43947 56797 43959 56831
rect 43901 56791 43959 56797
rect 43990 56788 43996 56840
rect 44048 56828 44054 56840
rect 44177 56831 44235 56837
rect 44177 56828 44189 56831
rect 44048 56800 44189 56828
rect 44048 56788 44054 56800
rect 44177 56797 44189 56800
rect 44223 56797 44235 56831
rect 45186 56828 45192 56840
rect 45147 56800 45192 56828
rect 44177 56791 44235 56797
rect 45186 56788 45192 56800
rect 45244 56788 45250 56840
rect 45922 56788 45928 56840
rect 45980 56828 45986 56840
rect 46017 56831 46075 56837
rect 46017 56828 46029 56831
rect 45980 56800 46029 56828
rect 45980 56788 45986 56800
rect 46017 56797 46029 56800
rect 46063 56797 46075 56831
rect 46017 56791 46075 56797
rect 48685 56831 48743 56837
rect 48685 56797 48697 56831
rect 48731 56797 48743 56831
rect 55490 56828 55496 56840
rect 55451 56800 55496 56828
rect 48685 56791 48743 56797
rect 39301 56763 39359 56769
rect 39301 56760 39313 56763
rect 38396 56732 39313 56760
rect 39301 56729 39313 56732
rect 39347 56760 39359 56763
rect 44358 56760 44364 56772
rect 39347 56732 44364 56760
rect 39347 56729 39359 56732
rect 39301 56723 39359 56729
rect 44358 56720 44364 56732
rect 44416 56720 44422 56772
rect 45370 56720 45376 56772
rect 45428 56760 45434 56772
rect 48700 56760 48728 56791
rect 55490 56788 55496 56800
rect 55548 56788 55554 56840
rect 45428 56732 48728 56760
rect 45428 56720 45434 56732
rect 39114 56692 39120 56704
rect 38304 56664 39120 56692
rect 39114 56652 39120 56664
rect 39172 56652 39178 56704
rect 40034 56692 40040 56704
rect 39995 56664 40040 56692
rect 40034 56652 40040 56664
rect 40092 56652 40098 56704
rect 40218 56652 40224 56704
rect 40276 56692 40282 56704
rect 41230 56692 41236 56704
rect 40276 56664 41236 56692
rect 40276 56652 40282 56664
rect 41230 56652 41236 56664
rect 41288 56652 41294 56704
rect 42886 56652 42892 56704
rect 42944 56692 42950 56704
rect 45833 56695 45891 56701
rect 45833 56692 45845 56695
rect 42944 56664 45845 56692
rect 42944 56652 42950 56664
rect 45833 56661 45845 56664
rect 45879 56661 45891 56695
rect 45833 56655 45891 56661
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 23198 56448 23204 56500
rect 23256 56488 23262 56500
rect 23385 56491 23443 56497
rect 23385 56488 23397 56491
rect 23256 56460 23397 56488
rect 23256 56448 23262 56460
rect 23385 56457 23397 56460
rect 23431 56457 23443 56491
rect 23385 56451 23443 56457
rect 23474 56448 23480 56500
rect 23532 56488 23538 56500
rect 26418 56488 26424 56500
rect 23532 56460 26424 56488
rect 23532 56448 23538 56460
rect 26418 56448 26424 56460
rect 26476 56488 26482 56500
rect 27154 56488 27160 56500
rect 26476 56460 27160 56488
rect 26476 56448 26482 56460
rect 27154 56448 27160 56460
rect 27212 56448 27218 56500
rect 27614 56488 27620 56500
rect 27575 56460 27620 56488
rect 27614 56448 27620 56460
rect 27672 56448 27678 56500
rect 27798 56448 27804 56500
rect 27856 56488 27862 56500
rect 28261 56491 28319 56497
rect 28261 56488 28273 56491
rect 27856 56460 28273 56488
rect 27856 56448 27862 56460
rect 28261 56457 28273 56460
rect 28307 56457 28319 56491
rect 28261 56451 28319 56457
rect 28994 56448 29000 56500
rect 29052 56488 29058 56500
rect 29089 56491 29147 56497
rect 29089 56488 29101 56491
rect 29052 56460 29101 56488
rect 29052 56448 29058 56460
rect 29089 56457 29101 56460
rect 29135 56457 29147 56491
rect 29089 56451 29147 56457
rect 30006 56448 30012 56500
rect 30064 56448 30070 56500
rect 30558 56448 30564 56500
rect 30616 56488 30622 56500
rect 30837 56491 30895 56497
rect 30837 56488 30849 56491
rect 30616 56460 30849 56488
rect 30616 56448 30622 56460
rect 30837 56457 30849 56460
rect 30883 56457 30895 56491
rect 30837 56451 30895 56457
rect 30926 56448 30932 56500
rect 30984 56488 30990 56500
rect 31938 56488 31944 56500
rect 30984 56460 31944 56488
rect 30984 56448 30990 56460
rect 31938 56448 31944 56460
rect 31996 56448 32002 56500
rect 32585 56491 32643 56497
rect 32585 56457 32597 56491
rect 32631 56488 32643 56491
rect 32950 56488 32956 56500
rect 32631 56460 32956 56488
rect 32631 56457 32643 56460
rect 32585 56451 32643 56457
rect 32950 56448 32956 56460
rect 33008 56448 33014 56500
rect 34146 56448 34152 56500
rect 34204 56448 34210 56500
rect 35342 56448 35348 56500
rect 35400 56488 35406 56500
rect 38746 56488 38752 56500
rect 35400 56460 38752 56488
rect 35400 56448 35406 56460
rect 38746 56448 38752 56460
rect 38804 56448 38810 56500
rect 42150 56488 42156 56500
rect 39132 56460 42156 56488
rect 25774 56420 25780 56432
rect 6886 56392 25780 56420
rect 5442 56312 5448 56364
rect 5500 56352 5506 56364
rect 6886 56352 6914 56392
rect 5500 56324 6914 56352
rect 5500 56312 5506 56324
rect 22554 56312 22560 56364
rect 22612 56352 22618 56364
rect 22649 56355 22707 56361
rect 22649 56352 22661 56355
rect 22612 56324 22661 56352
rect 22612 56312 22618 56324
rect 22649 56321 22661 56324
rect 22695 56321 22707 56355
rect 23566 56352 23572 56364
rect 23527 56324 23572 56352
rect 22649 56315 22707 56321
rect 23566 56312 23572 56324
rect 23624 56312 23630 56364
rect 23934 56312 23940 56364
rect 23992 56352 23998 56364
rect 24044 56361 24072 56392
rect 25774 56380 25780 56392
rect 25832 56420 25838 56432
rect 27632 56420 27660 56448
rect 25832 56392 26280 56420
rect 25832 56380 25838 56392
rect 24029 56355 24087 56361
rect 24029 56352 24041 56355
rect 23992 56324 24041 56352
rect 23992 56312 23998 56324
rect 24029 56321 24041 56324
rect 24075 56321 24087 56355
rect 24029 56315 24087 56321
rect 25409 56355 25467 56361
rect 25409 56321 25421 56355
rect 25455 56352 25467 56355
rect 25682 56352 25688 56364
rect 25455 56324 25688 56352
rect 25455 56321 25467 56324
rect 25409 56315 25467 56321
rect 25682 56312 25688 56324
rect 25740 56312 25746 56364
rect 26252 56361 26280 56392
rect 26436 56392 27660 56420
rect 26436 56361 26464 56392
rect 28350 56380 28356 56432
rect 28408 56420 28414 56432
rect 30024 56420 30052 56448
rect 31846 56420 31852 56432
rect 28408 56392 30052 56420
rect 31220 56392 31852 56420
rect 28408 56380 28414 56392
rect 26237 56355 26295 56361
rect 26237 56321 26249 56355
rect 26283 56321 26295 56355
rect 26237 56315 26295 56321
rect 26421 56355 26479 56361
rect 26421 56321 26433 56355
rect 26467 56321 26479 56355
rect 27246 56352 27252 56364
rect 26421 56315 26479 56321
rect 26528 56324 26924 56352
rect 27207 56324 27252 56352
rect 23658 56244 23664 56296
rect 23716 56284 23722 56296
rect 24305 56287 24363 56293
rect 24305 56284 24317 56287
rect 23716 56256 24317 56284
rect 23716 56244 23722 56256
rect 24305 56253 24317 56256
rect 24351 56284 24363 56287
rect 25222 56284 25228 56296
rect 24351 56256 25228 56284
rect 24351 56253 24363 56256
rect 24305 56247 24363 56253
rect 25222 56244 25228 56256
rect 25280 56244 25286 56296
rect 17126 56176 17132 56228
rect 17184 56216 17190 56228
rect 26528 56216 26556 56324
rect 26602 56244 26608 56296
rect 26660 56284 26666 56296
rect 26660 56256 26705 56284
rect 26660 56244 26666 56256
rect 17184 56188 26556 56216
rect 26896 56216 26924 56324
rect 27246 56312 27252 56324
rect 27304 56312 27310 56364
rect 27338 56312 27344 56364
rect 27396 56352 27402 56364
rect 27676 56355 27734 56361
rect 27676 56352 27688 56355
rect 27396 56324 27688 56352
rect 27396 56312 27402 56324
rect 27676 56321 27688 56324
rect 27722 56352 27734 56355
rect 28442 56352 28448 56364
rect 27722 56324 28304 56352
rect 28403 56324 28448 56352
rect 27722 56321 27734 56324
rect 27676 56315 27734 56321
rect 27154 56284 27160 56296
rect 27115 56256 27160 56284
rect 27154 56244 27160 56256
rect 27212 56244 27218 56296
rect 27801 56219 27859 56225
rect 27801 56216 27813 56219
rect 26896 56188 27813 56216
rect 17184 56176 17190 56188
rect 27801 56185 27813 56188
rect 27847 56185 27859 56219
rect 28276 56216 28304 56324
rect 28442 56312 28448 56324
rect 28500 56312 28506 56364
rect 28629 56355 28687 56361
rect 28629 56321 28641 56355
rect 28675 56352 28687 56355
rect 29089 56355 29147 56361
rect 29089 56352 29101 56355
rect 28675 56324 29101 56352
rect 28675 56321 28687 56324
rect 28629 56315 28687 56321
rect 29089 56321 29101 56324
rect 29135 56352 29147 56355
rect 29270 56352 29276 56364
rect 29135 56324 29276 56352
rect 29135 56321 29147 56324
rect 29089 56315 29147 56321
rect 29270 56312 29276 56324
rect 29328 56312 29334 56364
rect 29362 56312 29368 56364
rect 29420 56352 29426 56364
rect 29420 56324 29465 56352
rect 29420 56312 29426 56324
rect 29914 56312 29920 56364
rect 29972 56352 29978 56364
rect 31220 56361 31248 56392
rect 31846 56380 31852 56392
rect 31904 56420 31910 56432
rect 33226 56420 33232 56432
rect 31904 56392 33232 56420
rect 31904 56380 31910 56392
rect 33226 56380 33232 56392
rect 33284 56380 33290 56432
rect 34164 56420 34192 56448
rect 35526 56420 35532 56432
rect 33336 56392 34192 56420
rect 34624 56392 35532 56420
rect 30009 56355 30067 56361
rect 30009 56352 30021 56355
rect 29972 56324 30021 56352
rect 29972 56312 29978 56324
rect 30009 56321 30021 56324
rect 30055 56321 30067 56355
rect 30009 56315 30067 56321
rect 31205 56355 31263 56361
rect 31205 56321 31217 56355
rect 31251 56321 31263 56355
rect 31205 56315 31263 56321
rect 31297 56355 31355 56361
rect 31297 56321 31309 56355
rect 31343 56352 31355 56355
rect 32306 56352 32312 56364
rect 31343 56324 32312 56352
rect 31343 56321 31355 56324
rect 31297 56315 31355 56321
rect 32306 56312 32312 56324
rect 32364 56312 32370 56364
rect 32677 56355 32735 56361
rect 32677 56321 32689 56355
rect 32723 56352 32735 56355
rect 32766 56352 32772 56364
rect 32723 56324 32772 56352
rect 32723 56321 32735 56324
rect 32677 56315 32735 56321
rect 32766 56312 32772 56324
rect 32824 56312 32830 56364
rect 32858 56312 32864 56364
rect 32916 56352 32922 56364
rect 33336 56361 33364 56392
rect 33321 56355 33379 56361
rect 33321 56352 33333 56355
rect 32916 56324 33333 56352
rect 32916 56312 32922 56324
rect 33321 56321 33333 56324
rect 33367 56321 33379 56355
rect 33321 56315 33379 56321
rect 33413 56355 33471 56361
rect 33413 56321 33425 56355
rect 33459 56321 33471 56355
rect 33413 56315 33471 56321
rect 28460 56284 28488 56312
rect 29181 56287 29239 56293
rect 29181 56284 29193 56287
rect 28460 56256 29193 56284
rect 29181 56253 29193 56256
rect 29227 56253 29239 56287
rect 29181 56247 29239 56253
rect 30834 56244 30840 56296
rect 30892 56284 30898 56296
rect 31021 56287 31079 56293
rect 31021 56284 31033 56287
rect 30892 56256 31033 56284
rect 30892 56244 30898 56256
rect 31021 56253 31033 56256
rect 31067 56253 31079 56287
rect 31021 56247 31079 56253
rect 31110 56244 31116 56296
rect 31168 56284 31174 56296
rect 33428 56284 33456 56315
rect 33502 56312 33508 56364
rect 33560 56352 33566 56364
rect 33597 56355 33655 56361
rect 33597 56352 33609 56355
rect 33560 56324 33609 56352
rect 33560 56312 33566 56324
rect 33597 56321 33609 56324
rect 33643 56321 33655 56355
rect 33597 56315 33655 56321
rect 33689 56355 33747 56361
rect 33689 56321 33701 56355
rect 33735 56352 33747 56355
rect 34149 56355 34207 56361
rect 34149 56352 34161 56355
rect 33735 56324 34161 56352
rect 33735 56321 33747 56324
rect 33689 56315 33747 56321
rect 34149 56321 34161 56324
rect 34195 56321 34207 56355
rect 34330 56352 34336 56364
rect 34291 56324 34336 56352
rect 34149 56315 34207 56321
rect 34330 56312 34336 56324
rect 34388 56312 34394 56364
rect 34624 56361 34652 56392
rect 35526 56380 35532 56392
rect 35584 56420 35590 56432
rect 36262 56420 36268 56432
rect 35584 56392 36268 56420
rect 35584 56380 35590 56392
rect 36262 56380 36268 56392
rect 36320 56380 36326 56432
rect 36446 56420 36452 56432
rect 36407 56392 36452 56420
rect 36446 56380 36452 56392
rect 36504 56380 36510 56432
rect 36722 56380 36728 56432
rect 36780 56420 36786 56432
rect 36817 56423 36875 56429
rect 36817 56420 36829 56423
rect 36780 56392 36829 56420
rect 36780 56380 36786 56392
rect 36817 56389 36829 56392
rect 36863 56389 36875 56423
rect 36817 56383 36875 56389
rect 37734 56380 37740 56432
rect 37792 56420 37798 56432
rect 39132 56420 39160 56460
rect 42150 56448 42156 56460
rect 42208 56448 42214 56500
rect 42702 56448 42708 56500
rect 42760 56488 42766 56500
rect 43717 56491 43775 56497
rect 43717 56488 43729 56491
rect 42760 56460 43729 56488
rect 42760 56448 42766 56460
rect 43717 56457 43729 56460
rect 43763 56488 43775 56491
rect 43990 56488 43996 56500
rect 43763 56460 43996 56488
rect 43763 56457 43775 56460
rect 43717 56451 43775 56457
rect 43990 56448 43996 56460
rect 44048 56448 44054 56500
rect 45370 56488 45376 56500
rect 44192 56460 45376 56488
rect 37792 56392 39160 56420
rect 37792 56380 37798 56392
rect 39206 56380 39212 56432
rect 39264 56420 39270 56432
rect 39942 56420 39948 56432
rect 39264 56392 39948 56420
rect 39264 56380 39270 56392
rect 39942 56380 39948 56392
rect 40000 56380 40006 56432
rect 40034 56380 40040 56432
rect 40092 56420 40098 56432
rect 40313 56423 40371 56429
rect 40313 56420 40325 56423
rect 40092 56392 40325 56420
rect 40092 56380 40098 56392
rect 40313 56389 40325 56392
rect 40359 56389 40371 56423
rect 40313 56383 40371 56389
rect 40405 56423 40463 56429
rect 40405 56389 40417 56423
rect 40451 56420 40463 56423
rect 44085 56423 44143 56429
rect 44085 56420 44097 56423
rect 40451 56392 44097 56420
rect 40451 56389 40463 56392
rect 40405 56383 40463 56389
rect 44085 56389 44097 56392
rect 44131 56389 44143 56423
rect 44085 56383 44143 56389
rect 34609 56355 34667 56361
rect 34609 56321 34621 56355
rect 34655 56321 34667 56355
rect 35710 56352 35716 56364
rect 35671 56324 35716 56352
rect 34609 56315 34667 56321
rect 34624 56284 34652 56315
rect 35710 56312 35716 56324
rect 35768 56312 35774 56364
rect 35802 56312 35808 56364
rect 35860 56352 35866 56364
rect 35860 56324 35905 56352
rect 35860 56312 35866 56324
rect 36538 56312 36544 56364
rect 36596 56352 36602 56364
rect 36633 56355 36691 56361
rect 36633 56352 36645 56355
rect 36596 56324 36645 56352
rect 36596 56312 36602 56324
rect 36633 56321 36645 56324
rect 36679 56321 36691 56355
rect 36633 56315 36691 56321
rect 36906 56312 36912 56364
rect 36964 56352 36970 56364
rect 38841 56355 38899 56361
rect 36964 56324 37009 56352
rect 36964 56312 36970 56324
rect 38841 56321 38853 56355
rect 38887 56352 38899 56355
rect 38887 56324 39344 56352
rect 38887 56321 38899 56324
rect 38841 56315 38899 56321
rect 31168 56256 31213 56284
rect 33428 56256 34652 56284
rect 31168 56244 31174 56256
rect 34698 56244 34704 56296
rect 34756 56284 34762 56296
rect 35820 56284 35848 56312
rect 34756 56256 35848 56284
rect 38197 56287 38255 56293
rect 34756 56244 34762 56256
rect 38197 56253 38209 56287
rect 38243 56284 38255 56287
rect 38286 56284 38292 56296
rect 38243 56256 38292 56284
rect 38243 56253 38255 56256
rect 38197 56247 38255 56253
rect 38286 56244 38292 56256
rect 38344 56284 38350 56296
rect 38657 56287 38715 56293
rect 38657 56284 38669 56287
rect 38344 56256 38669 56284
rect 38344 56244 38350 56256
rect 38657 56253 38669 56256
rect 38703 56253 38715 56287
rect 38657 56247 38715 56253
rect 39025 56287 39083 56293
rect 39025 56253 39037 56287
rect 39071 56284 39083 56287
rect 39206 56284 39212 56296
rect 39071 56256 39212 56284
rect 39071 56253 39083 56256
rect 39025 56247 39083 56253
rect 39206 56244 39212 56256
rect 39264 56244 39270 56296
rect 31570 56216 31576 56228
rect 28276 56188 31576 56216
rect 27801 56179 27859 56185
rect 31570 56176 31576 56188
rect 31628 56176 31634 56228
rect 34054 56176 34060 56228
rect 34112 56216 34118 56228
rect 34790 56216 34796 56228
rect 34112 56188 34796 56216
rect 34112 56176 34118 56188
rect 34790 56176 34796 56188
rect 34848 56176 34854 56228
rect 34882 56176 34888 56228
rect 34940 56216 34946 56228
rect 35710 56216 35716 56228
rect 34940 56188 35716 56216
rect 34940 56176 34946 56188
rect 35710 56176 35716 56188
rect 35768 56176 35774 56228
rect 37921 56219 37979 56225
rect 37921 56185 37933 56219
rect 37967 56216 37979 56219
rect 39114 56216 39120 56228
rect 37967 56188 39120 56216
rect 37967 56185 37979 56188
rect 37921 56179 37979 56185
rect 39114 56176 39120 56188
rect 39172 56176 39178 56228
rect 39316 56216 39344 56324
rect 40126 56312 40132 56364
rect 40184 56361 40190 56364
rect 40184 56355 40233 56361
rect 40184 56321 40187 56355
rect 40221 56321 40233 56355
rect 40184 56315 40233 56321
rect 40184 56312 40190 56315
rect 40034 56284 40040 56296
rect 39995 56256 40040 56284
rect 40034 56244 40040 56256
rect 40092 56244 40098 56296
rect 40328 56284 40356 56383
rect 40494 56352 40500 56364
rect 40455 56324 40500 56352
rect 40494 56312 40500 56324
rect 40552 56312 40558 56364
rect 41601 56355 41659 56361
rect 40604 56324 41414 56352
rect 40604 56284 40632 56324
rect 40328 56256 40632 56284
rect 40681 56287 40739 56293
rect 40681 56253 40693 56287
rect 40727 56284 40739 56287
rect 40770 56284 40776 56296
rect 40727 56256 40776 56284
rect 40727 56253 40739 56256
rect 40681 56247 40739 56253
rect 40770 56244 40776 56256
rect 40828 56244 40834 56296
rect 41386 56284 41414 56324
rect 41601 56321 41613 56355
rect 41647 56352 41659 56355
rect 42613 56355 42671 56361
rect 42613 56352 42625 56355
rect 41647 56324 42625 56352
rect 41647 56321 41659 56324
rect 41601 56315 41659 56321
rect 42613 56321 42625 56324
rect 42659 56321 42671 56355
rect 42613 56315 42671 56321
rect 42702 56312 42708 56364
rect 42760 56352 42766 56364
rect 42797 56355 42855 56361
rect 42797 56352 42809 56355
rect 42760 56324 42809 56352
rect 42760 56312 42766 56324
rect 42797 56321 42809 56324
rect 42843 56321 42855 56355
rect 42797 56315 42855 56321
rect 42889 56355 42947 56361
rect 42889 56321 42901 56355
rect 42935 56321 42947 56355
rect 43070 56352 43076 56364
rect 43031 56324 43076 56352
rect 42889 56315 42947 56321
rect 41877 56287 41935 56293
rect 41877 56284 41889 56287
rect 41386 56256 41889 56284
rect 41877 56253 41889 56256
rect 41923 56284 41935 56287
rect 41966 56284 41972 56296
rect 41923 56256 41972 56284
rect 41923 56253 41935 56256
rect 41877 56247 41935 56253
rect 41966 56244 41972 56256
rect 42024 56284 42030 56296
rect 42426 56284 42432 56296
rect 42024 56256 42432 56284
rect 42024 56244 42030 56256
rect 42426 56244 42432 56256
rect 42484 56244 42490 56296
rect 42518 56244 42524 56296
rect 42576 56284 42582 56296
rect 42904 56284 42932 56315
rect 43070 56312 43076 56324
rect 43128 56312 43134 56364
rect 43162 56312 43168 56364
rect 43220 56352 43226 56364
rect 43622 56352 43628 56364
rect 43220 56324 43265 56352
rect 43583 56324 43628 56352
rect 43220 56312 43226 56324
rect 43622 56312 43628 56324
rect 43680 56312 43686 56364
rect 43898 56352 43904 56364
rect 43811 56324 43904 56352
rect 43898 56312 43904 56324
rect 43956 56352 43962 56364
rect 44192 56352 44220 56460
rect 45370 56448 45376 56460
rect 45428 56448 45434 56500
rect 49694 56448 49700 56500
rect 49752 56488 49758 56500
rect 50157 56491 50215 56497
rect 50157 56488 50169 56491
rect 49752 56460 50169 56488
rect 49752 56448 49758 56460
rect 50157 56457 50169 56460
rect 50203 56457 50215 56491
rect 51442 56488 51448 56500
rect 51403 56460 51448 56488
rect 50157 56451 50215 56457
rect 51442 56448 51448 56460
rect 51500 56448 51506 56500
rect 53006 56488 53012 56500
rect 52967 56460 53012 56488
rect 53006 56448 53012 56460
rect 53064 56448 53070 56500
rect 54754 56448 54760 56500
rect 54812 56488 54818 56500
rect 55490 56488 55496 56500
rect 54812 56460 55496 56488
rect 54812 56448 54818 56460
rect 55490 56448 55496 56460
rect 55548 56448 55554 56500
rect 45646 56420 45652 56432
rect 43956 56324 44220 56352
rect 44284 56392 45652 56420
rect 43956 56312 43962 56324
rect 43254 56284 43260 56296
rect 42576 56256 43260 56284
rect 42576 56244 42582 56256
rect 43254 56244 43260 56256
rect 43312 56284 43318 56296
rect 44284 56284 44312 56392
rect 45646 56380 45652 56392
rect 45704 56380 45710 56432
rect 44910 56352 44916 56364
rect 44871 56324 44916 56352
rect 44910 56312 44916 56324
rect 44968 56312 44974 56364
rect 45738 56312 45744 56364
rect 45796 56361 45802 56364
rect 45796 56355 45829 56361
rect 45817 56321 45829 56355
rect 45796 56315 45829 56321
rect 45925 56355 45983 56361
rect 45925 56321 45937 56355
rect 45971 56321 45983 56355
rect 45925 56315 45983 56321
rect 45796 56312 45802 56315
rect 44818 56284 44824 56296
rect 43312 56256 44312 56284
rect 44779 56256 44824 56284
rect 43312 56244 43318 56256
rect 44818 56244 44824 56256
rect 44876 56244 44882 56296
rect 45940 56284 45968 56315
rect 46474 56312 46480 56364
rect 46532 56352 46538 56364
rect 47029 56355 47087 56361
rect 47029 56352 47041 56355
rect 46532 56324 47041 56352
rect 46532 56312 46538 56324
rect 47029 56321 47041 56324
rect 47075 56321 47087 56355
rect 47029 56315 47087 56321
rect 47854 56312 47860 56364
rect 47912 56352 47918 56364
rect 47949 56355 48007 56361
rect 47949 56352 47961 56355
rect 47912 56324 47961 56352
rect 47912 56312 47918 56324
rect 47949 56321 47961 56324
rect 47995 56321 48007 56355
rect 47949 56315 48007 56321
rect 48774 56312 48780 56364
rect 48832 56352 48838 56364
rect 48869 56355 48927 56361
rect 48869 56352 48881 56355
rect 48832 56324 48881 56352
rect 48832 56312 48838 56324
rect 48869 56321 48881 56324
rect 48915 56321 48927 56355
rect 48869 56315 48927 56321
rect 49234 56312 49240 56364
rect 49292 56352 49298 56364
rect 49513 56355 49571 56361
rect 49513 56352 49525 56355
rect 49292 56324 49525 56352
rect 49292 56312 49298 56324
rect 49513 56321 49525 56324
rect 49559 56321 49571 56355
rect 49513 56315 49571 56321
rect 46842 56284 46848 56296
rect 45940 56256 46848 56284
rect 46842 56244 46848 56256
rect 46900 56244 46906 56296
rect 39390 56216 39396 56228
rect 39303 56188 39396 56216
rect 39390 56176 39396 56188
rect 39448 56216 39454 56228
rect 44545 56219 44603 56225
rect 44545 56216 44557 56219
rect 39448 56188 44557 56216
rect 39448 56176 39454 56188
rect 44545 56185 44557 56188
rect 44591 56185 44603 56219
rect 44545 56179 44603 56185
rect 44634 56176 44640 56228
rect 44692 56216 44698 56228
rect 46385 56219 46443 56225
rect 46385 56216 46397 56219
rect 44692 56188 46397 56216
rect 44692 56176 44698 56188
rect 46385 56185 46397 56188
rect 46431 56185 46443 56219
rect 46385 56179 46443 56185
rect 25498 56108 25504 56160
rect 25556 56148 25562 56160
rect 25593 56151 25651 56157
rect 25593 56148 25605 56151
rect 25556 56120 25605 56148
rect 25556 56108 25562 56120
rect 25593 56117 25605 56120
rect 25639 56117 25651 56151
rect 25593 56111 25651 56117
rect 25682 56108 25688 56160
rect 25740 56148 25746 56160
rect 32490 56148 32496 56160
rect 25740 56120 32496 56148
rect 25740 56108 25746 56120
rect 32490 56108 32496 56120
rect 32548 56108 32554 56160
rect 33134 56148 33140 56160
rect 33095 56120 33140 56148
rect 33134 56108 33140 56120
rect 33192 56108 33198 56160
rect 33594 56108 33600 56160
rect 33652 56148 33658 56160
rect 34422 56148 34428 56160
rect 33652 56120 34428 56148
rect 33652 56108 33658 56120
rect 34422 56108 34428 56120
rect 34480 56108 34486 56160
rect 34517 56151 34575 56157
rect 34517 56117 34529 56151
rect 34563 56148 34575 56151
rect 34900 56148 34928 56176
rect 35618 56148 35624 56160
rect 34563 56120 34928 56148
rect 35579 56120 35624 56148
rect 34563 56117 34575 56120
rect 34517 56111 34575 56117
rect 35618 56108 35624 56120
rect 35676 56108 35682 56160
rect 36814 56108 36820 56160
rect 36872 56148 36878 56160
rect 37737 56151 37795 56157
rect 37737 56148 37749 56151
rect 36872 56120 37749 56148
rect 36872 56108 36878 56120
rect 37737 56117 37749 56120
rect 37783 56117 37795 56151
rect 37737 56111 37795 56117
rect 37826 56108 37832 56160
rect 37884 56148 37890 56160
rect 39577 56151 39635 56157
rect 39577 56148 39589 56151
rect 37884 56120 39589 56148
rect 37884 56108 37890 56120
rect 39577 56117 39589 56120
rect 39623 56148 39635 56151
rect 40954 56148 40960 56160
rect 39623 56120 40960 56148
rect 39623 56117 39635 56120
rect 39577 56111 39635 56117
rect 40954 56108 40960 56120
rect 41012 56108 41018 56160
rect 41414 56108 41420 56160
rect 41472 56148 41478 56160
rect 41782 56148 41788 56160
rect 41472 56120 41517 56148
rect 41743 56120 41788 56148
rect 41472 56108 41478 56120
rect 41782 56108 41788 56120
rect 41840 56108 41846 56160
rect 43070 56108 43076 56160
rect 43128 56148 43134 56160
rect 45462 56148 45468 56160
rect 43128 56120 45468 56148
rect 43128 56108 43134 56120
rect 45462 56108 45468 56120
rect 45520 56108 45526 56160
rect 45738 56148 45744 56160
rect 45699 56120 45744 56148
rect 45738 56108 45744 56120
rect 45796 56108 45802 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 23750 55904 23756 55956
rect 23808 55944 23814 55956
rect 23845 55947 23903 55953
rect 23845 55944 23857 55947
rect 23808 55916 23857 55944
rect 23808 55904 23814 55916
rect 23845 55913 23857 55916
rect 23891 55913 23903 55947
rect 23845 55907 23903 55913
rect 24673 55947 24731 55953
rect 24673 55913 24685 55947
rect 24719 55944 24731 55947
rect 25038 55944 25044 55956
rect 24719 55916 25044 55944
rect 24719 55913 24731 55916
rect 24673 55907 24731 55913
rect 25038 55904 25044 55916
rect 25096 55904 25102 55956
rect 27985 55947 28043 55953
rect 27985 55913 27997 55947
rect 28031 55944 28043 55947
rect 28442 55944 28448 55956
rect 28031 55916 28448 55944
rect 28031 55913 28043 55916
rect 27985 55907 28043 55913
rect 28442 55904 28448 55916
rect 28500 55904 28506 55956
rect 30374 55944 30380 55956
rect 28552 55916 30380 55944
rect 28552 55876 28580 55916
rect 30374 55904 30380 55916
rect 30432 55904 30438 55956
rect 31570 55944 31576 55956
rect 31531 55916 31576 55944
rect 31570 55904 31576 55916
rect 31628 55904 31634 55956
rect 34333 55947 34391 55953
rect 34333 55944 34345 55947
rect 31726 55916 34345 55944
rect 31726 55876 31754 55916
rect 34333 55913 34345 55916
rect 34379 55913 34391 55947
rect 34333 55907 34391 55913
rect 34422 55904 34428 55956
rect 34480 55944 34486 55956
rect 35897 55947 35955 55953
rect 35897 55944 35909 55947
rect 34480 55916 35909 55944
rect 34480 55904 34486 55916
rect 35897 55913 35909 55916
rect 35943 55913 35955 55947
rect 35897 55907 35955 55913
rect 36906 55904 36912 55956
rect 36964 55944 36970 55956
rect 37001 55947 37059 55953
rect 37001 55944 37013 55947
rect 36964 55916 37013 55944
rect 36964 55904 36970 55916
rect 37001 55913 37013 55916
rect 37047 55913 37059 55947
rect 37001 55907 37059 55913
rect 37645 55947 37703 55953
rect 37645 55913 37657 55947
rect 37691 55944 37703 55947
rect 37826 55944 37832 55956
rect 37691 55916 37832 55944
rect 37691 55913 37703 55916
rect 37645 55907 37703 55913
rect 37826 55904 37832 55916
rect 37884 55904 37890 55956
rect 39025 55947 39083 55953
rect 39025 55913 39037 55947
rect 39071 55944 39083 55947
rect 39114 55944 39120 55956
rect 39071 55916 39120 55944
rect 39071 55913 39083 55916
rect 39025 55907 39083 55913
rect 39114 55904 39120 55916
rect 39172 55904 39178 55956
rect 40037 55947 40095 55953
rect 40037 55913 40049 55947
rect 40083 55944 40095 55947
rect 40126 55944 40132 55956
rect 40083 55916 40132 55944
rect 40083 55913 40095 55916
rect 40037 55907 40095 55913
rect 40126 55904 40132 55916
rect 40184 55904 40190 55956
rect 40494 55904 40500 55956
rect 40552 55944 40558 55956
rect 41601 55947 41659 55953
rect 41601 55944 41613 55947
rect 40552 55916 41613 55944
rect 40552 55904 40558 55916
rect 41601 55913 41613 55916
rect 41647 55913 41659 55947
rect 41601 55907 41659 55913
rect 41874 55904 41880 55956
rect 41932 55944 41938 55956
rect 42613 55947 42671 55953
rect 42613 55944 42625 55947
rect 41932 55916 42625 55944
rect 41932 55904 41938 55916
rect 42613 55913 42625 55916
rect 42659 55944 42671 55947
rect 42702 55944 42708 55956
rect 42659 55916 42708 55944
rect 42659 55913 42671 55916
rect 42613 55907 42671 55913
rect 42702 55904 42708 55916
rect 42760 55904 42766 55956
rect 42981 55947 43039 55953
rect 42981 55913 42993 55947
rect 43027 55944 43039 55947
rect 43162 55944 43168 55956
rect 43027 55916 43168 55944
rect 43027 55913 43039 55916
rect 42981 55907 43039 55913
rect 43162 55904 43168 55916
rect 43220 55904 43226 55956
rect 43438 55944 43444 55956
rect 43399 55916 43444 55944
rect 43438 55904 43444 55916
rect 43496 55904 43502 55956
rect 46842 55944 46848 55956
rect 46803 55916 46848 55944
rect 46842 55904 46848 55916
rect 46900 55904 46906 55956
rect 26712 55848 28580 55876
rect 28644 55848 31754 55876
rect 31864 55848 32352 55876
rect 23385 55811 23443 55817
rect 23385 55777 23397 55811
rect 23431 55808 23443 55811
rect 25222 55808 25228 55820
rect 23431 55780 25228 55808
rect 23431 55777 23443 55780
rect 23385 55771 23443 55777
rect 25222 55768 25228 55780
rect 25280 55808 25286 55820
rect 25685 55811 25743 55817
rect 25685 55808 25697 55811
rect 25280 55780 25697 55808
rect 25280 55768 25286 55780
rect 25685 55777 25697 55780
rect 25731 55808 25743 55811
rect 26237 55811 26295 55817
rect 26237 55808 26249 55811
rect 25731 55780 26249 55808
rect 25731 55777 25743 55780
rect 25685 55771 25743 55777
rect 26237 55777 26249 55780
rect 26283 55808 26295 55811
rect 26510 55808 26516 55820
rect 26283 55780 26516 55808
rect 26283 55777 26295 55780
rect 26237 55771 26295 55777
rect 26510 55768 26516 55780
rect 26568 55808 26574 55820
rect 26712 55817 26740 55848
rect 28644 55817 28672 55848
rect 26697 55811 26755 55817
rect 26697 55808 26709 55811
rect 26568 55780 26709 55808
rect 26568 55768 26574 55780
rect 26697 55777 26709 55780
rect 26743 55777 26755 55811
rect 28629 55811 28687 55817
rect 28629 55808 28641 55811
rect 26697 55771 26755 55777
rect 28000 55780 28641 55808
rect 24026 55740 24032 55752
rect 23987 55712 24032 55740
rect 24026 55700 24032 55712
rect 24084 55700 24090 55752
rect 24857 55743 24915 55749
rect 24857 55709 24869 55743
rect 24903 55740 24915 55743
rect 25317 55743 25375 55749
rect 25317 55740 25329 55743
rect 24903 55712 25329 55740
rect 24903 55709 24915 55712
rect 24857 55703 24915 55709
rect 25317 55709 25329 55712
rect 25363 55709 25375 55743
rect 25317 55703 25375 55709
rect 25501 55743 25559 55749
rect 25501 55709 25513 55743
rect 25547 55740 25559 55743
rect 25590 55740 25596 55752
rect 25547 55712 25596 55740
rect 25547 55709 25559 55712
rect 25501 55703 25559 55709
rect 25590 55700 25596 55712
rect 25648 55700 25654 55752
rect 26881 55743 26939 55749
rect 26881 55709 26893 55743
rect 26927 55740 26939 55743
rect 27338 55740 27344 55752
rect 26927 55712 27344 55740
rect 26927 55709 26939 55712
rect 26881 55703 26939 55709
rect 27338 55700 27344 55712
rect 27396 55700 27402 55752
rect 28000 55749 28028 55780
rect 28629 55777 28641 55780
rect 28675 55777 28687 55811
rect 28629 55771 28687 55777
rect 28721 55811 28779 55817
rect 28721 55777 28733 55811
rect 28767 55808 28779 55811
rect 29917 55811 29975 55817
rect 29917 55808 29929 55811
rect 28767 55780 29929 55808
rect 28767 55777 28779 55780
rect 28721 55771 28779 55777
rect 29917 55777 29929 55780
rect 29963 55777 29975 55811
rect 29917 55771 29975 55777
rect 27709 55743 27767 55749
rect 27709 55709 27721 55743
rect 27755 55709 27767 55743
rect 27709 55703 27767 55709
rect 27985 55743 28043 55749
rect 27985 55709 27997 55743
rect 28031 55709 28043 55743
rect 27985 55703 28043 55709
rect 27065 55607 27123 55613
rect 27065 55573 27077 55607
rect 27111 55604 27123 55607
rect 27154 55604 27160 55616
rect 27111 55576 27160 55604
rect 27111 55573 27123 55576
rect 27065 55567 27123 55573
rect 27154 55564 27160 55576
rect 27212 55564 27218 55616
rect 27724 55604 27752 55703
rect 28350 55700 28356 55752
rect 28408 55740 28414 55752
rect 28537 55743 28595 55749
rect 28537 55740 28549 55743
rect 28408 55712 28549 55740
rect 28408 55700 28414 55712
rect 28537 55709 28549 55712
rect 28583 55709 28595 55743
rect 28537 55703 28595 55709
rect 27801 55675 27859 55681
rect 27801 55641 27813 55675
rect 27847 55672 27859 55675
rect 28442 55672 28448 55684
rect 27847 55644 28448 55672
rect 27847 55641 27859 55644
rect 27801 55635 27859 55641
rect 28442 55632 28448 55644
rect 28500 55672 28506 55684
rect 28736 55672 28764 55771
rect 30006 55768 30012 55820
rect 30064 55808 30070 55820
rect 30742 55808 30748 55820
rect 30064 55780 30748 55808
rect 30064 55768 30070 55780
rect 30742 55768 30748 55780
rect 30800 55808 30806 55820
rect 31110 55808 31116 55820
rect 30800 55780 31116 55808
rect 30800 55768 30806 55780
rect 31110 55768 31116 55780
rect 31168 55808 31174 55820
rect 31864 55808 31892 55848
rect 31168 55780 31892 55808
rect 32324 55808 32352 55848
rect 32490 55836 32496 55888
rect 32548 55876 32554 55888
rect 32953 55879 33011 55885
rect 32953 55876 32965 55879
rect 32548 55848 32965 55876
rect 32548 55836 32554 55848
rect 32953 55845 32965 55848
rect 32999 55845 33011 55879
rect 34698 55876 34704 55888
rect 32953 55839 33011 55845
rect 33428 55848 34704 55876
rect 32766 55808 32772 55820
rect 32324 55780 32772 55808
rect 31168 55768 31174 55780
rect 28813 55743 28871 55749
rect 28813 55709 28825 55743
rect 28859 55740 28871 55743
rect 28994 55740 29000 55752
rect 28859 55712 29000 55740
rect 28859 55709 28871 55712
rect 28813 55703 28871 55709
rect 28500 55644 28764 55672
rect 28500 55632 28506 55644
rect 28828 55604 28856 55703
rect 28994 55700 29000 55712
rect 29052 55700 29058 55752
rect 30926 55740 30932 55752
rect 30887 55712 30932 55740
rect 30926 55700 30932 55712
rect 30984 55700 30990 55752
rect 31220 55749 31248 55780
rect 32766 55768 32772 55780
rect 32824 55808 32830 55820
rect 33428 55817 33456 55848
rect 34698 55836 34704 55848
rect 34756 55836 34762 55888
rect 34882 55876 34888 55888
rect 34843 55848 34888 55876
rect 34882 55836 34888 55848
rect 34940 55836 34946 55888
rect 38194 55836 38200 55888
rect 38252 55876 38258 55888
rect 40865 55879 40923 55885
rect 40865 55876 40877 55879
rect 38252 55848 40877 55876
rect 38252 55836 38258 55848
rect 40865 55845 40877 55848
rect 40911 55845 40923 55879
rect 40865 55839 40923 55845
rect 40954 55836 40960 55888
rect 41012 55876 41018 55888
rect 41012 55848 41414 55876
rect 41012 55836 41018 55848
rect 33413 55811 33471 55817
rect 33413 55808 33425 55811
rect 32824 55780 33425 55808
rect 32824 55768 32830 55780
rect 33413 55777 33425 55780
rect 33459 55777 33471 55811
rect 35158 55808 35164 55820
rect 35119 55780 35164 55808
rect 33413 55771 33471 55777
rect 35158 55768 35164 55780
rect 35216 55768 35222 55820
rect 36814 55808 36820 55820
rect 36775 55780 36820 55808
rect 36814 55768 36820 55780
rect 36872 55768 36878 55820
rect 41386 55808 41414 55848
rect 44358 55836 44364 55888
rect 44416 55876 44422 55888
rect 45462 55876 45468 55888
rect 44416 55848 44461 55876
rect 45423 55848 45468 55876
rect 44416 55836 44422 55848
rect 45462 55836 45468 55848
rect 45520 55836 45526 55888
rect 45557 55879 45615 55885
rect 45557 55845 45569 55879
rect 45603 55876 45615 55879
rect 45646 55876 45652 55888
rect 45603 55848 45652 55876
rect 45603 55845 45615 55848
rect 45557 55839 45615 55845
rect 45646 55836 45652 55848
rect 45704 55836 45710 55888
rect 51810 55808 51816 55820
rect 41386 55780 51816 55808
rect 51810 55768 51816 55780
rect 51868 55768 51874 55820
rect 31205 55743 31263 55749
rect 31205 55709 31217 55743
rect 31251 55709 31263 55743
rect 31386 55740 31392 55752
rect 31347 55712 31392 55740
rect 31205 55703 31263 55709
rect 31386 55700 31392 55712
rect 31444 55700 31450 55752
rect 32217 55743 32275 55749
rect 32217 55709 32229 55743
rect 32263 55709 32275 55743
rect 32217 55703 32275 55709
rect 32493 55743 32551 55749
rect 32493 55709 32505 55743
rect 32539 55740 32551 55743
rect 32582 55740 32588 55752
rect 32539 55712 32588 55740
rect 32539 55709 32551 55712
rect 32493 55703 32551 55709
rect 30098 55672 30104 55684
rect 30059 55644 30104 55672
rect 30098 55632 30104 55644
rect 30156 55632 30162 55684
rect 30282 55672 30288 55684
rect 30243 55644 30288 55672
rect 30282 55632 30288 55644
rect 30340 55632 30346 55684
rect 31018 55632 31024 55684
rect 31076 55681 31082 55684
rect 31076 55675 31125 55681
rect 31076 55641 31079 55675
rect 31113 55641 31125 55675
rect 31076 55635 31125 55641
rect 31297 55675 31355 55681
rect 31297 55641 31309 55675
rect 31343 55672 31355 55675
rect 32033 55675 32091 55681
rect 32033 55672 32045 55675
rect 31343 55644 32045 55672
rect 31343 55641 31355 55644
rect 31297 55635 31355 55641
rect 32033 55641 32045 55644
rect 32079 55641 32091 55675
rect 32033 55635 32091 55641
rect 31076 55632 31082 55635
rect 27724 55576 28856 55604
rect 28997 55607 29055 55613
rect 28997 55573 29009 55607
rect 29043 55604 29055 55607
rect 29270 55604 29276 55616
rect 29043 55576 29276 55604
rect 29043 55573 29055 55576
rect 28997 55567 29055 55573
rect 29270 55564 29276 55576
rect 29328 55564 29334 55616
rect 30006 55564 30012 55616
rect 30064 55604 30070 55616
rect 30300 55604 30328 55632
rect 30064 55576 30328 55604
rect 32232 55604 32260 55703
rect 32582 55700 32588 55712
rect 32640 55700 32646 55752
rect 33134 55740 33140 55752
rect 33095 55712 33140 55740
rect 33134 55700 33140 55712
rect 33192 55700 33198 55752
rect 33226 55700 33232 55752
rect 33284 55740 33290 55752
rect 33321 55743 33379 55749
rect 33321 55740 33333 55743
rect 33284 55712 33333 55740
rect 33284 55700 33290 55712
rect 33321 55709 33333 55712
rect 33367 55709 33379 55743
rect 34054 55740 34060 55752
rect 34015 55712 34060 55740
rect 33321 55703 33379 55709
rect 34054 55700 34060 55712
rect 34112 55700 34118 55752
rect 34149 55743 34207 55749
rect 34149 55709 34161 55743
rect 34195 55740 34207 55743
rect 34238 55740 34244 55752
rect 34195 55712 34244 55740
rect 34195 55709 34207 55712
rect 34149 55703 34207 55709
rect 34238 55700 34244 55712
rect 34296 55700 34302 55752
rect 34422 55750 34428 55752
rect 34351 55749 34428 55750
rect 34333 55743 34428 55749
rect 34333 55709 34345 55743
rect 34379 55722 34428 55743
rect 34379 55709 34391 55722
rect 34333 55703 34391 55709
rect 34422 55700 34428 55722
rect 34480 55700 34486 55752
rect 34606 55700 34612 55752
rect 34664 55740 34670 55752
rect 35253 55743 35311 55749
rect 35253 55740 35265 55743
rect 34664 55712 35265 55740
rect 34664 55700 34670 55712
rect 35253 55709 35265 55712
rect 35299 55709 35311 55743
rect 35253 55703 35311 55709
rect 36725 55743 36783 55749
rect 36725 55709 36737 55743
rect 36771 55740 36783 55743
rect 38105 55743 38163 55749
rect 38105 55740 38117 55743
rect 36771 55712 38117 55740
rect 36771 55709 36783 55712
rect 36725 55703 36783 55709
rect 38105 55709 38117 55712
rect 38151 55709 38163 55743
rect 38105 55703 38163 55709
rect 38194 55700 38200 55752
rect 38252 55740 38258 55752
rect 38289 55743 38347 55749
rect 38289 55740 38301 55743
rect 38252 55712 38301 55740
rect 38252 55700 38258 55712
rect 38289 55709 38301 55712
rect 38335 55709 38347 55743
rect 38562 55740 38568 55752
rect 38475 55712 38568 55740
rect 38289 55703 38347 55709
rect 38562 55700 38568 55712
rect 38620 55740 38626 55752
rect 42518 55740 42524 55752
rect 38620 55712 40448 55740
rect 42479 55712 42524 55740
rect 38620 55700 38626 55712
rect 40420 55684 40448 55712
rect 42518 55700 42524 55712
rect 42576 55700 42582 55752
rect 42797 55743 42855 55749
rect 42797 55709 42809 55743
rect 42843 55740 42855 55743
rect 42886 55740 42892 55752
rect 42843 55712 42892 55740
rect 42843 55709 42855 55712
rect 42797 55703 42855 55709
rect 42886 55700 42892 55712
rect 42944 55700 42950 55752
rect 43990 55700 43996 55752
rect 44048 55740 44054 55752
rect 44085 55743 44143 55749
rect 44085 55740 44097 55743
rect 44048 55712 44097 55740
rect 44048 55700 44054 55712
rect 44085 55709 44097 55712
rect 44131 55740 44143 55743
rect 44361 55743 44419 55749
rect 44131 55712 44220 55740
rect 44131 55709 44143 55712
rect 44085 55703 44143 55709
rect 32398 55632 32404 55684
rect 32456 55672 32462 55684
rect 32858 55672 32864 55684
rect 32456 55644 32864 55672
rect 32456 55632 32462 55644
rect 32858 55632 32864 55644
rect 32916 55632 32922 55684
rect 39209 55675 39267 55681
rect 39209 55641 39221 55675
rect 39255 55641 39267 55675
rect 39390 55672 39396 55684
rect 39351 55644 39396 55672
rect 39209 55635 39267 55641
rect 35342 55604 35348 55616
rect 32232 55576 35348 55604
rect 30064 55564 30070 55576
rect 35342 55564 35348 55576
rect 35400 55564 35406 55616
rect 38470 55604 38476 55616
rect 38431 55576 38476 55604
rect 38470 55564 38476 55576
rect 38528 55564 38534 55616
rect 39224 55604 39252 55635
rect 39390 55632 39396 55644
rect 39448 55632 39454 55684
rect 40218 55672 40224 55684
rect 40179 55644 40224 55672
rect 40218 55632 40224 55644
rect 40276 55632 40282 55684
rect 40402 55672 40408 55684
rect 40363 55644 40408 55672
rect 40402 55632 40408 55644
rect 40460 55632 40466 55684
rect 41785 55675 41843 55681
rect 41785 55641 41797 55675
rect 41831 55672 41843 55675
rect 41874 55672 41880 55684
rect 41831 55644 41880 55672
rect 41831 55641 41843 55644
rect 41785 55635 41843 55641
rect 41874 55632 41880 55644
rect 41932 55632 41938 55684
rect 41969 55675 42027 55681
rect 41969 55641 41981 55675
rect 42015 55672 42027 55675
rect 43622 55672 43628 55684
rect 42015 55644 43628 55672
rect 42015 55641 42027 55644
rect 41969 55635 42027 55641
rect 39298 55604 39304 55616
rect 39224 55576 39304 55604
rect 39298 55564 39304 55576
rect 39356 55564 39362 55616
rect 39482 55564 39488 55616
rect 39540 55604 39546 55616
rect 41984 55604 42012 55635
rect 43622 55632 43628 55644
rect 43680 55632 43686 55684
rect 44192 55672 44220 55712
rect 44361 55709 44373 55743
rect 44407 55740 44419 55743
rect 44818 55740 44824 55752
rect 44407 55712 44824 55740
rect 44407 55709 44419 55712
rect 44361 55703 44419 55709
rect 44818 55700 44824 55712
rect 44876 55740 44882 55752
rect 45189 55743 45247 55749
rect 45189 55740 45201 55743
rect 44876 55712 45201 55740
rect 44876 55700 44882 55712
rect 45189 55709 45201 55712
rect 45235 55709 45247 55743
rect 45370 55740 45376 55752
rect 45331 55712 45376 55740
rect 45189 55703 45247 55709
rect 45370 55700 45376 55712
rect 45428 55700 45434 55752
rect 45649 55743 45707 55749
rect 45649 55709 45661 55743
rect 45695 55709 45707 55743
rect 45649 55703 45707 55709
rect 45664 55672 45692 55703
rect 45738 55672 45744 55684
rect 44192 55644 45744 55672
rect 45738 55632 45744 55644
rect 45796 55632 45802 55684
rect 39540 55576 42012 55604
rect 44177 55607 44235 55613
rect 39540 55564 39546 55576
rect 44177 55573 44189 55607
rect 44223 55604 44235 55607
rect 44910 55604 44916 55616
rect 44223 55576 44916 55604
rect 44223 55573 44235 55576
rect 44177 55567 44235 55573
rect 44910 55564 44916 55576
rect 44968 55564 44974 55616
rect 46198 55604 46204 55616
rect 46159 55576 46204 55604
rect 46198 55564 46204 55576
rect 46256 55564 46262 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 23934 55400 23940 55412
rect 23895 55372 23940 55400
rect 23934 55360 23940 55372
rect 23992 55360 23998 55412
rect 25130 55360 25136 55412
rect 25188 55400 25194 55412
rect 25685 55403 25743 55409
rect 25685 55400 25697 55403
rect 25188 55372 25697 55400
rect 25188 55360 25194 55372
rect 25685 55369 25697 55372
rect 25731 55369 25743 55403
rect 26418 55400 26424 55412
rect 26379 55372 26424 55400
rect 25685 55363 25743 55369
rect 26418 55360 26424 55372
rect 26476 55360 26482 55412
rect 27246 55360 27252 55412
rect 27304 55400 27310 55412
rect 27341 55403 27399 55409
rect 27341 55400 27353 55403
rect 27304 55372 27353 55400
rect 27304 55360 27310 55372
rect 27341 55369 27353 55372
rect 27387 55369 27399 55403
rect 27341 55363 27399 55369
rect 27985 55403 28043 55409
rect 27985 55369 27997 55403
rect 28031 55400 28043 55403
rect 30834 55400 30840 55412
rect 28031 55372 30840 55400
rect 28031 55369 28043 55372
rect 27985 55363 28043 55369
rect 30834 55360 30840 55372
rect 30892 55360 30898 55412
rect 30929 55403 30987 55409
rect 30929 55369 30941 55403
rect 30975 55400 30987 55403
rect 31018 55400 31024 55412
rect 30975 55372 31024 55400
rect 30975 55369 30987 55372
rect 30929 55363 30987 55369
rect 31018 55360 31024 55372
rect 31076 55360 31082 55412
rect 31386 55360 31392 55412
rect 31444 55400 31450 55412
rect 32309 55403 32367 55409
rect 32309 55400 32321 55403
rect 31444 55372 32321 55400
rect 31444 55360 31450 55372
rect 32309 55369 32321 55372
rect 32355 55369 32367 55403
rect 32309 55363 32367 55369
rect 32674 55360 32680 55412
rect 32732 55400 32738 55412
rect 33778 55400 33784 55412
rect 32732 55372 33784 55400
rect 32732 55360 32738 55372
rect 33778 55360 33784 55372
rect 33836 55360 33842 55412
rect 33962 55360 33968 55412
rect 34020 55400 34026 55412
rect 34425 55403 34483 55409
rect 34425 55400 34437 55403
rect 34020 55372 34437 55400
rect 34020 55360 34026 55372
rect 34425 55369 34437 55372
rect 34471 55369 34483 55403
rect 34425 55363 34483 55369
rect 34606 55360 34612 55412
rect 34664 55400 34670 55412
rect 35069 55403 35127 55409
rect 35069 55400 35081 55403
rect 34664 55372 35081 55400
rect 34664 55360 34670 55372
rect 35069 55369 35081 55372
rect 35115 55400 35127 55403
rect 35158 55400 35164 55412
rect 35115 55372 35164 55400
rect 35115 55369 35127 55372
rect 35069 55363 35127 55369
rect 35158 55360 35164 55372
rect 35216 55360 35222 55412
rect 36630 55400 36636 55412
rect 35268 55372 36636 55400
rect 24489 55335 24547 55341
rect 24489 55301 24501 55335
rect 24535 55332 24547 55335
rect 25041 55335 25099 55341
rect 25041 55332 25053 55335
rect 24535 55304 25053 55332
rect 24535 55301 24547 55304
rect 24489 55295 24547 55301
rect 25041 55301 25053 55304
rect 25087 55332 25099 55335
rect 25222 55332 25228 55344
rect 25087 55304 25228 55332
rect 25087 55301 25099 55304
rect 25041 55295 25099 55301
rect 25222 55292 25228 55304
rect 25280 55292 25286 55344
rect 29089 55335 29147 55341
rect 29089 55301 29101 55335
rect 29135 55332 29147 55335
rect 29730 55332 29736 55344
rect 29135 55304 29736 55332
rect 29135 55301 29147 55304
rect 29089 55295 29147 55301
rect 29730 55292 29736 55304
rect 29788 55292 29794 55344
rect 30098 55292 30104 55344
rect 30156 55332 30162 55344
rect 33980 55332 34008 55360
rect 30156 55304 32812 55332
rect 30156 55292 30162 55304
rect 25498 55264 25504 55276
rect 25459 55236 25504 55264
rect 25498 55224 25504 55236
rect 25556 55224 25562 55276
rect 26602 55264 26608 55276
rect 26563 55236 26608 55264
rect 26602 55224 26608 55236
rect 26660 55224 26666 55276
rect 27154 55264 27160 55276
rect 27115 55236 27160 55264
rect 27154 55224 27160 55236
rect 27212 55224 27218 55276
rect 27798 55264 27804 55276
rect 27711 55236 27804 55264
rect 27798 55224 27804 55236
rect 27856 55264 27862 55276
rect 28902 55264 28908 55276
rect 27856 55236 28908 55264
rect 27856 55224 27862 55236
rect 28902 55224 28908 55236
rect 28960 55224 28966 55276
rect 29270 55264 29276 55276
rect 29231 55236 29276 55264
rect 29270 55224 29276 55236
rect 29328 55224 29334 55276
rect 29365 55267 29423 55273
rect 29365 55233 29377 55267
rect 29411 55264 29423 55267
rect 30006 55264 30012 55276
rect 29411 55236 29868 55264
rect 29967 55236 30012 55264
rect 29411 55233 29423 55236
rect 29365 55227 29423 55233
rect 28629 55199 28687 55205
rect 28629 55165 28641 55199
rect 28675 55196 28687 55199
rect 29454 55196 29460 55208
rect 28675 55168 29460 55196
rect 28675 55165 28687 55168
rect 28629 55159 28687 55165
rect 29454 55156 29460 55168
rect 29512 55156 29518 55208
rect 29840 55196 29868 55236
rect 30006 55224 30012 55236
rect 30064 55224 30070 55276
rect 30208 55273 30236 55304
rect 30193 55267 30251 55273
rect 30193 55233 30205 55267
rect 30239 55233 30251 55267
rect 30193 55227 30251 55233
rect 31018 55224 31024 55276
rect 31076 55264 31082 55276
rect 31113 55267 31171 55273
rect 31113 55264 31125 55267
rect 31076 55236 31125 55264
rect 31076 55224 31082 55236
rect 31113 55233 31125 55236
rect 31159 55233 31171 55267
rect 31113 55227 31171 55233
rect 31202 55224 31208 55276
rect 31260 55264 31266 55276
rect 31297 55267 31355 55273
rect 31297 55264 31309 55267
rect 31260 55236 31309 55264
rect 31260 55224 31266 55236
rect 31297 55233 31309 55236
rect 31343 55233 31355 55267
rect 31297 55227 31355 55233
rect 32398 55224 32404 55276
rect 32456 55264 32462 55276
rect 32493 55267 32551 55273
rect 32493 55264 32505 55267
rect 32456 55236 32505 55264
rect 32456 55224 32462 55236
rect 32493 55233 32505 55236
rect 32539 55233 32551 55267
rect 32674 55264 32680 55276
rect 32635 55236 32680 55264
rect 32493 55227 32551 55233
rect 32674 55224 32680 55236
rect 32732 55224 32738 55276
rect 32784 55264 32812 55304
rect 33060 55304 34008 55332
rect 33060 55264 33088 55304
rect 32784 55236 33088 55264
rect 33318 55224 33324 55276
rect 33376 55264 33382 55276
rect 34514 55264 34520 55276
rect 33376 55236 34520 55264
rect 33376 55224 33382 55236
rect 34514 55224 34520 55236
rect 34572 55264 34578 55276
rect 35268 55273 35296 55372
rect 36630 55360 36636 55372
rect 36688 55360 36694 55412
rect 38470 55360 38476 55412
rect 38528 55400 38534 55412
rect 38528 55372 38654 55400
rect 38528 55360 38534 55372
rect 35434 55292 35440 55344
rect 35492 55332 35498 55344
rect 38626 55332 38654 55372
rect 40034 55360 40040 55412
rect 40092 55400 40098 55412
rect 40135 55403 40193 55409
rect 40135 55400 40147 55403
rect 40092 55372 40147 55400
rect 40092 55360 40098 55372
rect 40135 55369 40147 55372
rect 40181 55369 40193 55403
rect 42794 55400 42800 55412
rect 40135 55363 40193 55369
rect 41386 55372 42800 55400
rect 39209 55335 39267 55341
rect 39209 55332 39221 55335
rect 35492 55304 36124 55332
rect 38626 55304 39221 55332
rect 35492 55292 35498 55304
rect 34609 55267 34667 55273
rect 34609 55264 34621 55267
rect 34572 55236 34621 55264
rect 34572 55224 34578 55236
rect 34609 55233 34621 55236
rect 34655 55233 34667 55267
rect 34609 55227 34667 55233
rect 35253 55267 35311 55273
rect 35253 55233 35265 55267
rect 35299 55264 35311 55267
rect 35342 55264 35348 55276
rect 35299 55236 35348 55264
rect 35299 55233 35311 55236
rect 35253 55227 35311 55233
rect 35342 55224 35348 55236
rect 35400 55224 35406 55276
rect 35529 55267 35587 55273
rect 35529 55233 35541 55267
rect 35575 55264 35587 55267
rect 35618 55264 35624 55276
rect 35575 55236 35624 55264
rect 35575 55233 35587 55236
rect 35529 55227 35587 55233
rect 35618 55224 35624 55236
rect 35676 55224 35682 55276
rect 31220 55196 31248 55224
rect 33778 55196 33784 55208
rect 29840 55168 31248 55196
rect 33739 55168 33784 55196
rect 33778 55156 33784 55168
rect 33836 55156 33842 55208
rect 36096 55205 36124 55304
rect 39209 55301 39221 55304
rect 39255 55301 39267 55335
rect 39209 55295 39267 55301
rect 39298 55292 39304 55344
rect 39356 55332 39362 55344
rect 41386 55332 41414 55372
rect 42794 55360 42800 55372
rect 42852 55360 42858 55412
rect 42886 55360 42892 55412
rect 42944 55400 42950 55412
rect 43990 55400 43996 55412
rect 42944 55372 43996 55400
rect 42944 55360 42950 55372
rect 43990 55360 43996 55372
rect 44048 55360 44054 55412
rect 44266 55400 44272 55412
rect 44227 55372 44272 55400
rect 44266 55360 44272 55372
rect 44324 55360 44330 55412
rect 45554 55360 45560 55412
rect 45612 55400 45618 55412
rect 46201 55403 46259 55409
rect 46201 55400 46213 55403
rect 45612 55372 46213 55400
rect 45612 55360 45618 55372
rect 46201 55369 46213 55372
rect 46247 55369 46259 55403
rect 46201 55363 46259 55369
rect 39356 55304 41414 55332
rect 39356 55292 39362 55304
rect 42334 55292 42340 55344
rect 42392 55332 42398 55344
rect 42392 55304 43668 55332
rect 42392 55292 42398 55304
rect 36998 55224 37004 55276
rect 37056 55264 37062 55276
rect 38194 55264 38200 55276
rect 37056 55236 37504 55264
rect 38155 55236 38200 55264
rect 37056 55224 37062 55236
rect 36081 55199 36139 55205
rect 36081 55165 36093 55199
rect 36127 55165 36139 55199
rect 36081 55159 36139 55165
rect 36354 55156 36360 55208
rect 36412 55196 36418 55208
rect 37476 55205 37504 55236
rect 38194 55224 38200 55236
rect 38252 55224 38258 55276
rect 38286 55224 38292 55276
rect 38344 55264 38350 55276
rect 38470 55264 38476 55276
rect 38344 55236 38389 55264
rect 38431 55236 38476 55264
rect 38344 55224 38350 55236
rect 38470 55224 38476 55236
rect 38528 55224 38534 55276
rect 38562 55224 38568 55276
rect 38620 55264 38626 55276
rect 39390 55264 39396 55276
rect 38620 55236 38665 55264
rect 39351 55236 39396 55264
rect 38620 55224 38626 55236
rect 39390 55224 39396 55236
rect 39448 55224 39454 55276
rect 39482 55224 39488 55276
rect 39540 55264 39546 55276
rect 39577 55267 39635 55273
rect 39577 55264 39589 55267
rect 39540 55236 39589 55264
rect 39540 55224 39546 55236
rect 39577 55233 39589 55236
rect 39623 55233 39635 55267
rect 39577 55227 39635 55233
rect 40037 55267 40095 55273
rect 40037 55233 40049 55267
rect 40083 55233 40095 55267
rect 40218 55264 40224 55276
rect 40179 55236 40224 55264
rect 40037 55227 40095 55233
rect 36725 55199 36783 55205
rect 36725 55196 36737 55199
rect 36412 55168 36737 55196
rect 36412 55156 36418 55168
rect 36725 55165 36737 55168
rect 36771 55165 36783 55199
rect 36725 55159 36783 55165
rect 37461 55199 37519 55205
rect 37461 55165 37473 55199
rect 37507 55165 37519 55199
rect 37461 55159 37519 55165
rect 38654 55156 38660 55208
rect 38712 55196 38718 55208
rect 38749 55199 38807 55205
rect 38749 55196 38761 55199
rect 38712 55168 38761 55196
rect 38712 55156 38718 55168
rect 38749 55165 38761 55168
rect 38795 55165 38807 55199
rect 38749 55159 38807 55165
rect 39942 55156 39948 55208
rect 40000 55196 40006 55208
rect 40052 55196 40080 55227
rect 40218 55224 40224 55236
rect 40276 55224 40282 55276
rect 40313 55267 40371 55273
rect 40313 55233 40325 55267
rect 40359 55264 40371 55267
rect 40402 55264 40408 55276
rect 40359 55236 40408 55264
rect 40359 55233 40371 55236
rect 40313 55227 40371 55233
rect 40402 55224 40408 55236
rect 40460 55264 40466 55276
rect 41690 55264 41696 55276
rect 40460 55236 41696 55264
rect 40460 55224 40466 55236
rect 41690 55224 41696 55236
rect 41748 55224 41754 55276
rect 41785 55267 41843 55273
rect 41785 55233 41797 55267
rect 41831 55264 41843 55267
rect 42150 55264 42156 55276
rect 41831 55236 42156 55264
rect 41831 55233 41843 55236
rect 41785 55227 41843 55233
rect 42150 55224 42156 55236
rect 42208 55224 42214 55276
rect 42886 55264 42892 55276
rect 42847 55236 42892 55264
rect 42886 55224 42892 55236
rect 42944 55224 42950 55276
rect 42981 55267 43039 55273
rect 42981 55233 42993 55267
rect 43027 55233 43039 55267
rect 42981 55227 43039 55233
rect 43109 55267 43167 55273
rect 43109 55233 43121 55267
rect 43155 55264 43167 55267
rect 43254 55264 43260 55276
rect 43155 55236 43260 55264
rect 43155 55233 43167 55236
rect 43109 55227 43167 55233
rect 40773 55199 40831 55205
rect 40773 55196 40785 55199
rect 40000 55168 40785 55196
rect 40000 55156 40006 55168
rect 40773 55165 40785 55168
rect 40819 55165 40831 55199
rect 40773 55159 40831 55165
rect 32214 55088 32220 55140
rect 32272 55128 32278 55140
rect 33137 55131 33195 55137
rect 33137 55128 33149 55131
rect 32272 55100 33149 55128
rect 32272 55088 32278 55100
rect 33137 55097 33149 55100
rect 33183 55097 33195 55131
rect 33137 55091 33195 55097
rect 35345 55131 35403 55137
rect 35345 55097 35357 55131
rect 35391 55097 35403 55131
rect 35345 55091 35403 55097
rect 35437 55131 35495 55137
rect 35437 55097 35449 55131
rect 35483 55128 35495 55131
rect 35526 55128 35532 55140
rect 35483 55100 35532 55128
rect 35483 55097 35495 55100
rect 35437 55091 35495 55097
rect 29086 55060 29092 55072
rect 29047 55032 29092 55060
rect 29086 55020 29092 55032
rect 29144 55020 29150 55072
rect 29822 55060 29828 55072
rect 29783 55032 29828 55060
rect 29822 55020 29828 55032
rect 29880 55020 29886 55072
rect 34698 55020 34704 55072
rect 34756 55060 34762 55072
rect 35360 55060 35388 55091
rect 35526 55088 35532 55100
rect 35584 55088 35590 55140
rect 37366 55088 37372 55140
rect 37424 55128 37430 55140
rect 42996 55128 43024 55227
rect 43254 55224 43260 55236
rect 43312 55224 43318 55276
rect 43640 55273 43668 55304
rect 44082 55292 44088 55344
rect 44140 55332 44146 55344
rect 45741 55335 45799 55341
rect 44140 55304 45692 55332
rect 44140 55292 44146 55304
rect 43625 55267 43683 55273
rect 43625 55233 43637 55267
rect 43671 55233 43683 55267
rect 43625 55227 43683 55233
rect 44174 55224 44180 55276
rect 44232 55264 44238 55276
rect 44453 55267 44511 55273
rect 44453 55264 44465 55267
rect 44232 55236 44465 55264
rect 44232 55224 44238 55236
rect 44453 55233 44465 55236
rect 44499 55264 44511 55267
rect 44913 55267 44971 55273
rect 44913 55264 44925 55267
rect 44499 55236 44925 55264
rect 44499 55233 44511 55236
rect 44453 55227 44511 55233
rect 44913 55233 44925 55236
rect 44959 55233 44971 55267
rect 45664 55264 45692 55304
rect 45741 55301 45753 55335
rect 45787 55332 45799 55335
rect 45922 55332 45928 55344
rect 45787 55304 45928 55332
rect 45787 55301 45799 55304
rect 45741 55295 45799 55301
rect 45922 55292 45928 55304
rect 45980 55292 45986 55344
rect 46198 55264 46204 55276
rect 45664 55236 46204 55264
rect 44913 55227 44971 55233
rect 46198 55224 46204 55236
rect 46256 55224 46262 55276
rect 53098 55196 53104 55208
rect 51046 55168 53104 55196
rect 43070 55128 43076 55140
rect 37424 55100 42932 55128
rect 42996 55100 43076 55128
rect 37424 55088 37430 55100
rect 34756 55032 35388 55060
rect 34756 55020 34762 55032
rect 41138 55020 41144 55072
rect 41196 55060 41202 55072
rect 41325 55063 41383 55069
rect 41325 55060 41337 55063
rect 41196 55032 41337 55060
rect 41196 55020 41202 55032
rect 41325 55029 41337 55032
rect 41371 55029 41383 55063
rect 41325 55023 41383 55029
rect 41693 55063 41751 55069
rect 41693 55029 41705 55063
rect 41739 55060 41751 55063
rect 42058 55060 42064 55072
rect 41739 55032 42064 55060
rect 41739 55029 41751 55032
rect 41693 55023 41751 55029
rect 42058 55020 42064 55032
rect 42116 55020 42122 55072
rect 42702 55060 42708 55072
rect 42663 55032 42708 55060
rect 42702 55020 42708 55032
rect 42760 55020 42766 55072
rect 42904 55060 42932 55100
rect 43070 55088 43076 55100
rect 43128 55088 43134 55140
rect 51046 55060 51074 55168
rect 53098 55156 53104 55168
rect 53156 55156 53162 55208
rect 42904 55032 51074 55060
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 25133 54859 25191 54865
rect 25133 54825 25145 54859
rect 25179 54856 25191 54859
rect 25222 54856 25228 54868
rect 25179 54828 25228 54856
rect 25179 54825 25191 54828
rect 25133 54819 25191 54825
rect 25222 54816 25228 54828
rect 25280 54816 25286 54868
rect 25774 54856 25780 54868
rect 25735 54828 25780 54856
rect 25774 54816 25780 54828
rect 25832 54816 25838 54868
rect 26513 54859 26571 54865
rect 26513 54825 26525 54859
rect 26559 54856 26571 54859
rect 26694 54856 26700 54868
rect 26559 54828 26700 54856
rect 26559 54825 26571 54828
rect 26513 54819 26571 54825
rect 26694 54816 26700 54828
rect 26752 54816 26758 54868
rect 27893 54859 27951 54865
rect 27893 54825 27905 54859
rect 27939 54856 27951 54859
rect 28074 54856 28080 54868
rect 27939 54828 28080 54856
rect 27939 54825 27951 54828
rect 27893 54819 27951 54825
rect 28074 54816 28080 54828
rect 28132 54816 28138 54868
rect 28994 54816 29000 54868
rect 29052 54856 29058 54868
rect 30285 54859 30343 54865
rect 30285 54856 30297 54859
rect 29052 54828 30297 54856
rect 29052 54816 29058 54828
rect 30285 54825 30297 54828
rect 30331 54825 30343 54859
rect 30285 54819 30343 54825
rect 30837 54859 30895 54865
rect 30837 54825 30849 54859
rect 30883 54856 30895 54859
rect 30926 54856 30932 54868
rect 30883 54828 30932 54856
rect 30883 54825 30895 54828
rect 30837 54819 30895 54825
rect 30926 54816 30932 54828
rect 30984 54816 30990 54868
rect 31938 54856 31944 54868
rect 31899 54828 31944 54856
rect 31938 54816 31944 54828
rect 31996 54816 32002 54868
rect 32122 54816 32128 54868
rect 32180 54856 32186 54868
rect 32861 54859 32919 54865
rect 32861 54856 32873 54859
rect 32180 54828 32873 54856
rect 32180 54816 32186 54828
rect 32861 54825 32873 54828
rect 32907 54856 32919 54859
rect 33597 54859 33655 54865
rect 33597 54856 33609 54859
rect 32907 54828 33609 54856
rect 32907 54825 32919 54828
rect 32861 54819 32919 54825
rect 33597 54825 33609 54828
rect 33643 54825 33655 54859
rect 33778 54856 33784 54868
rect 33739 54828 33784 54856
rect 33597 54819 33655 54825
rect 33778 54816 33784 54828
rect 33836 54816 33842 54868
rect 34790 54816 34796 54868
rect 34848 54856 34854 54868
rect 34885 54859 34943 54865
rect 34885 54856 34897 54859
rect 34848 54828 34897 54856
rect 34848 54816 34854 54828
rect 34885 54825 34897 54828
rect 34931 54825 34943 54859
rect 34885 54819 34943 54825
rect 35621 54859 35679 54865
rect 35621 54825 35633 54859
rect 35667 54856 35679 54859
rect 35802 54856 35808 54868
rect 35667 54828 35808 54856
rect 35667 54825 35679 54828
rect 35621 54819 35679 54825
rect 35802 54816 35808 54828
rect 35860 54856 35866 54868
rect 36173 54859 36231 54865
rect 36173 54856 36185 54859
rect 35860 54828 36185 54856
rect 35860 54816 35866 54828
rect 36173 54825 36185 54828
rect 36219 54856 36231 54859
rect 37277 54859 37335 54865
rect 37277 54856 37289 54859
rect 36219 54828 37289 54856
rect 36219 54825 36231 54828
rect 36173 54819 36231 54825
rect 37277 54825 37289 54828
rect 37323 54856 37335 54859
rect 37366 54856 37372 54868
rect 37323 54828 37372 54856
rect 37323 54825 37335 54828
rect 37277 54819 37335 54825
rect 37366 54816 37372 54828
rect 37424 54816 37430 54868
rect 38105 54859 38163 54865
rect 38105 54825 38117 54859
rect 38151 54856 38163 54859
rect 38194 54856 38200 54868
rect 38151 54828 38200 54856
rect 38151 54825 38163 54828
rect 38105 54819 38163 54825
rect 38194 54816 38200 54828
rect 38252 54816 38258 54868
rect 39485 54859 39543 54865
rect 39485 54825 39497 54859
rect 39531 54856 39543 54859
rect 40218 54856 40224 54868
rect 39531 54828 40224 54856
rect 39531 54825 39543 54828
rect 39485 54819 39543 54825
rect 40218 54816 40224 54828
rect 40276 54816 40282 54868
rect 40494 54816 40500 54868
rect 40552 54856 40558 54868
rect 40865 54859 40923 54865
rect 40865 54856 40877 54859
rect 40552 54828 40877 54856
rect 40552 54816 40558 54828
rect 40865 54825 40877 54828
rect 40911 54856 40923 54859
rect 41230 54856 41236 54868
rect 40911 54828 41236 54856
rect 40911 54825 40923 54828
rect 40865 54819 40923 54825
rect 41230 54816 41236 54828
rect 41288 54816 41294 54868
rect 41690 54856 41696 54868
rect 41651 54828 41696 54856
rect 41690 54816 41696 54828
rect 41748 54816 41754 54868
rect 28442 54788 28448 54800
rect 28403 54760 28448 54788
rect 28442 54748 28448 54760
rect 28500 54748 28506 54800
rect 35710 54748 35716 54800
rect 35768 54788 35774 54800
rect 36446 54788 36452 54800
rect 35768 54760 36452 54788
rect 35768 54748 35774 54760
rect 36446 54748 36452 54760
rect 36504 54788 36510 54800
rect 36725 54791 36783 54797
rect 36725 54788 36737 54791
rect 36504 54760 36737 54788
rect 36504 54748 36510 54760
rect 36725 54757 36737 54760
rect 36771 54788 36783 54791
rect 37826 54788 37832 54800
rect 36771 54760 37832 54788
rect 36771 54757 36783 54760
rect 36725 54751 36783 54757
rect 37826 54748 37832 54760
rect 37884 54748 37890 54800
rect 40034 54788 40040 54800
rect 39995 54760 40040 54788
rect 40034 54748 40040 54760
rect 40092 54748 40098 54800
rect 43717 54791 43775 54797
rect 43717 54788 43729 54791
rect 40144 54760 43729 54788
rect 28813 54723 28871 54729
rect 28813 54689 28825 54723
rect 28859 54720 28871 54723
rect 39209 54723 39267 54729
rect 39209 54720 39221 54723
rect 28859 54692 29868 54720
rect 28859 54689 28871 54692
rect 28813 54683 28871 54689
rect 29840 54664 29868 54692
rect 30116 54692 31156 54720
rect 25774 54612 25780 54664
rect 25832 54652 25838 54664
rect 26973 54655 27031 54661
rect 26973 54652 26985 54655
rect 25832 54624 26985 54652
rect 25832 54612 25838 54624
rect 26973 54621 26985 54624
rect 27019 54652 27031 54655
rect 27154 54652 27160 54664
rect 27019 54624 27160 54652
rect 27019 54621 27031 54624
rect 26973 54615 27031 54621
rect 27154 54612 27160 54624
rect 27212 54612 27218 54664
rect 29730 54652 29736 54664
rect 29691 54624 29736 54652
rect 29730 54612 29736 54624
rect 29788 54612 29794 54664
rect 29822 54612 29828 54664
rect 29880 54652 29886 54664
rect 30116 54661 30144 54692
rect 31128 54664 31156 54692
rect 38304 54692 39221 54720
rect 30009 54655 30067 54661
rect 29880 54624 29925 54652
rect 29880 54612 29886 54624
rect 30009 54621 30021 54655
rect 30055 54621 30067 54655
rect 30009 54615 30067 54621
rect 30101 54655 30159 54661
rect 30101 54621 30113 54655
rect 30147 54621 30159 54655
rect 30101 54615 30159 54621
rect 27065 54587 27123 54593
rect 27065 54553 27077 54587
rect 27111 54584 27123 54587
rect 27111 54556 28672 54584
rect 27111 54553 27123 54556
rect 27065 54547 27123 54553
rect 28353 54519 28411 54525
rect 28353 54485 28365 54519
rect 28399 54516 28411 54519
rect 28534 54516 28540 54528
rect 28399 54488 28540 54516
rect 28399 54485 28411 54488
rect 28353 54479 28411 54485
rect 28534 54476 28540 54488
rect 28592 54476 28598 54528
rect 28644 54516 28672 54556
rect 29270 54544 29276 54596
rect 29328 54584 29334 54596
rect 30024 54584 30052 54615
rect 30742 54612 30748 54664
rect 30800 54652 30806 54664
rect 30837 54655 30895 54661
rect 30837 54652 30849 54655
rect 30800 54624 30849 54652
rect 30800 54612 30806 54624
rect 30837 54621 30849 54624
rect 30883 54621 30895 54655
rect 31018 54652 31024 54664
rect 30979 54624 31024 54652
rect 30837 54615 30895 54621
rect 31018 54612 31024 54624
rect 31076 54612 31082 54664
rect 31110 54612 31116 54664
rect 31168 54652 31174 54664
rect 31757 54655 31815 54661
rect 31168 54624 31213 54652
rect 31168 54612 31174 54624
rect 31757 54621 31769 54655
rect 31803 54652 31815 54655
rect 31846 54652 31852 54664
rect 31803 54624 31852 54652
rect 31803 54621 31815 54624
rect 31757 54615 31815 54621
rect 31846 54612 31852 54624
rect 31904 54652 31910 54664
rect 32582 54652 32588 54664
rect 31904 54624 32588 54652
rect 31904 54612 31910 54624
rect 32582 54612 32588 54624
rect 32640 54612 32646 54664
rect 33134 54652 33140 54664
rect 33095 54624 33140 54652
rect 33134 54612 33140 54624
rect 33192 54612 33198 54664
rect 38304 54661 38332 54692
rect 39209 54689 39221 54692
rect 39255 54720 39267 54723
rect 39482 54720 39488 54732
rect 39255 54692 39488 54720
rect 39255 54689 39267 54692
rect 39209 54683 39267 54689
rect 39482 54680 39488 54692
rect 39540 54720 39546 54732
rect 40144 54720 40172 54760
rect 43717 54757 43729 54760
rect 43763 54757 43775 54791
rect 43717 54751 43775 54757
rect 41230 54720 41236 54732
rect 39540 54692 40172 54720
rect 41143 54692 41236 54720
rect 39540 54680 39546 54692
rect 41230 54680 41236 54692
rect 41288 54720 41294 54732
rect 42794 54720 42800 54732
rect 41288 54692 42196 54720
rect 42755 54692 42800 54720
rect 41288 54680 41294 54692
rect 38289 54655 38347 54661
rect 38289 54621 38301 54655
rect 38335 54621 38347 54655
rect 38289 54615 38347 54621
rect 38473 54655 38531 54661
rect 38473 54621 38485 54655
rect 38519 54652 38531 54655
rect 39117 54655 39175 54661
rect 39117 54652 39129 54655
rect 38519 54624 39129 54652
rect 38519 54621 38531 54624
rect 38473 54615 38531 54621
rect 39117 54621 39129 54624
rect 39163 54652 39175 54655
rect 39390 54652 39396 54664
rect 39163 54624 39396 54652
rect 39163 54621 39175 54624
rect 39117 54615 39175 54621
rect 39390 54612 39396 54624
rect 39448 54612 39454 54664
rect 40773 54655 40831 54661
rect 40773 54621 40785 54655
rect 40819 54652 40831 54655
rect 41877 54655 41935 54661
rect 40819 54624 41414 54652
rect 40819 54621 40831 54624
rect 40773 54615 40831 54621
rect 29328 54556 30052 54584
rect 29328 54544 29334 54556
rect 33318 54544 33324 54596
rect 33376 54584 33382 54596
rect 33749 54587 33807 54593
rect 33749 54584 33761 54587
rect 33376 54556 33761 54584
rect 33376 54544 33382 54556
rect 33749 54553 33761 54556
rect 33795 54553 33807 54587
rect 33962 54584 33968 54596
rect 33875 54556 33968 54584
rect 33749 54547 33807 54553
rect 33962 54544 33968 54556
rect 34020 54584 34026 54596
rect 34330 54584 34336 54596
rect 34020 54556 34336 54584
rect 34020 54544 34026 54556
rect 34330 54544 34336 54556
rect 34388 54544 34394 54596
rect 41386 54584 41414 54624
rect 41877 54621 41889 54655
rect 41923 54652 41935 54655
rect 42058 54652 42064 54664
rect 41923 54624 42064 54652
rect 41923 54621 41935 54624
rect 41877 54615 41935 54621
rect 42058 54612 42064 54624
rect 42116 54612 42122 54664
rect 42168 54661 42196 54692
rect 42794 54680 42800 54692
rect 42852 54680 42858 54732
rect 42889 54723 42947 54729
rect 42889 54689 42901 54723
rect 42935 54720 42947 54723
rect 43070 54720 43076 54732
rect 42935 54692 43076 54720
rect 42935 54689 42947 54692
rect 42889 54683 42947 54689
rect 42153 54655 42211 54661
rect 42153 54621 42165 54655
rect 42199 54621 42211 54655
rect 42153 54615 42211 54621
rect 42904 54584 42932 54683
rect 43070 54680 43076 54692
rect 43128 54680 43134 54732
rect 43254 54720 43260 54732
rect 43215 54692 43260 54720
rect 43254 54680 43260 54692
rect 43312 54680 43318 54732
rect 44174 54720 44180 54732
rect 44135 54692 44180 54720
rect 44174 54680 44180 54692
rect 44232 54680 44238 54732
rect 43898 54612 43904 54664
rect 43956 54652 43962 54664
rect 44085 54655 44143 54661
rect 44085 54652 44097 54655
rect 43956 54624 44097 54652
rect 43956 54612 43962 54624
rect 44085 54621 44097 54624
rect 44131 54621 44143 54655
rect 44085 54615 44143 54621
rect 41386 54556 42932 54584
rect 29362 54516 29368 54528
rect 28644 54488 29368 54516
rect 29362 54476 29368 54488
rect 29420 54476 29426 54528
rect 32214 54516 32220 54528
rect 32175 54488 32220 54516
rect 32214 54476 32220 54488
rect 32272 54476 32278 54528
rect 32490 54476 32496 54528
rect 32548 54516 32554 54528
rect 32677 54519 32735 54525
rect 32677 54516 32689 54519
rect 32548 54488 32689 54516
rect 32548 54476 32554 54488
rect 32677 54485 32689 54488
rect 32723 54485 32735 54519
rect 32677 54479 32735 54485
rect 42061 54519 42119 54525
rect 42061 54485 42073 54519
rect 42107 54516 42119 54519
rect 42150 54516 42156 54528
rect 42107 54488 42156 54516
rect 42107 54485 42119 54488
rect 42061 54479 42119 54485
rect 42150 54476 42156 54488
rect 42208 54476 42214 54528
rect 42610 54516 42616 54528
rect 42571 54488 42616 54516
rect 42610 54476 42616 54488
rect 42668 54476 42674 54528
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 26510 54312 26516 54324
rect 26471 54284 26516 54312
rect 26510 54272 26516 54284
rect 26568 54272 26574 54324
rect 27154 54312 27160 54324
rect 27115 54284 27160 54312
rect 27154 54272 27160 54284
rect 27212 54272 27218 54324
rect 27798 54312 27804 54324
rect 27759 54284 27804 54312
rect 27798 54272 27804 54284
rect 27856 54272 27862 54324
rect 28258 54312 28264 54324
rect 28219 54284 28264 54312
rect 28258 54272 28264 54284
rect 28316 54272 28322 54324
rect 29270 54272 29276 54324
rect 29328 54312 29334 54324
rect 29365 54315 29423 54321
rect 29365 54312 29377 54315
rect 29328 54284 29377 54312
rect 29328 54272 29334 54284
rect 29365 54281 29377 54284
rect 29411 54281 29423 54315
rect 29365 54275 29423 54281
rect 30742 54272 30748 54324
rect 30800 54312 30806 54324
rect 31205 54315 31263 54321
rect 31205 54312 31217 54315
rect 30800 54284 31217 54312
rect 30800 54272 30806 54284
rect 31205 54281 31217 54284
rect 31251 54281 31263 54315
rect 31205 54275 31263 54281
rect 32861 54315 32919 54321
rect 32861 54281 32873 54315
rect 32907 54312 32919 54315
rect 33226 54312 33232 54324
rect 32907 54284 33232 54312
rect 32907 54281 32919 54284
rect 32861 54275 32919 54281
rect 33226 54272 33232 54284
rect 33284 54272 33290 54324
rect 34330 54312 34336 54324
rect 34243 54284 34336 54312
rect 34330 54272 34336 54284
rect 34388 54312 34394 54324
rect 35526 54312 35532 54324
rect 34388 54284 35532 54312
rect 34388 54272 34394 54284
rect 35526 54272 35532 54284
rect 35584 54272 35590 54324
rect 36446 54312 36452 54324
rect 36407 54284 36452 54312
rect 36446 54272 36452 54284
rect 36504 54272 36510 54324
rect 37274 54272 37280 54324
rect 37332 54312 37338 54324
rect 37461 54315 37519 54321
rect 37461 54312 37473 54315
rect 37332 54284 37473 54312
rect 37332 54272 37338 54284
rect 37461 54281 37473 54284
rect 37507 54281 37519 54315
rect 37461 54275 37519 54281
rect 38930 54272 38936 54324
rect 38988 54312 38994 54324
rect 39117 54315 39175 54321
rect 39117 54312 39129 54315
rect 38988 54284 39129 54312
rect 38988 54272 38994 54284
rect 39117 54281 39129 54284
rect 39163 54281 39175 54315
rect 40494 54312 40500 54324
rect 40455 54284 40500 54312
rect 39117 54275 39175 54281
rect 40494 54272 40500 54284
rect 40552 54272 40558 54324
rect 41509 54315 41567 54321
rect 41509 54281 41521 54315
rect 41555 54312 41567 54315
rect 41782 54312 41788 54324
rect 41555 54284 41788 54312
rect 41555 54281 41567 54284
rect 41509 54275 41567 54281
rect 41782 54272 41788 54284
rect 41840 54272 41846 54324
rect 41966 54312 41972 54324
rect 41927 54284 41972 54312
rect 41966 54272 41972 54284
rect 42024 54272 42030 54324
rect 42702 54312 42708 54324
rect 42663 54284 42708 54312
rect 42702 54272 42708 54284
rect 42760 54272 42766 54324
rect 44174 54312 44180 54324
rect 44135 54284 44180 54312
rect 44174 54272 44180 54284
rect 44232 54272 44238 54324
rect 29549 54247 29607 54253
rect 29549 54213 29561 54247
rect 29595 54244 29607 54247
rect 32674 54244 32680 54256
rect 29595 54216 32680 54244
rect 29595 54213 29607 54216
rect 29549 54207 29607 54213
rect 28629 54179 28687 54185
rect 28629 54145 28641 54179
rect 28675 54176 28687 54179
rect 29086 54176 29092 54188
rect 28675 54148 29092 54176
rect 28675 54145 28687 54148
rect 28629 54139 28687 54145
rect 29086 54136 29092 54148
rect 29144 54136 29150 54188
rect 29733 54179 29791 54185
rect 29733 54145 29745 54179
rect 29779 54145 29791 54179
rect 29733 54139 29791 54145
rect 28534 54108 28540 54120
rect 28495 54080 28540 54108
rect 28534 54068 28540 54080
rect 28592 54068 28598 54120
rect 29748 54108 29776 54139
rect 30282 54136 30288 54188
rect 30340 54176 30346 54188
rect 30392 54185 30420 54216
rect 32674 54204 32680 54216
rect 32732 54204 32738 54256
rect 34514 54204 34520 54256
rect 34572 54244 34578 54256
rect 35897 54247 35955 54253
rect 35897 54244 35909 54247
rect 34572 54216 35909 54244
rect 34572 54204 34578 54216
rect 35897 54213 35909 54216
rect 35943 54213 35955 54247
rect 35897 54207 35955 54213
rect 42150 54204 42156 54256
rect 42208 54244 42214 54256
rect 43073 54247 43131 54253
rect 43073 54244 43085 54247
rect 42208 54216 43085 54244
rect 42208 54204 42214 54216
rect 43073 54213 43085 54216
rect 43119 54213 43131 54247
rect 43073 54207 43131 54213
rect 30377 54179 30435 54185
rect 30377 54176 30389 54179
rect 30340 54148 30389 54176
rect 30340 54136 30346 54148
rect 30377 54145 30389 54148
rect 30423 54145 30435 54179
rect 32490 54176 32496 54188
rect 32451 54148 32496 54176
rect 30377 54139 30435 54145
rect 32490 54136 32496 54148
rect 32548 54136 32554 54188
rect 33873 54179 33931 54185
rect 33873 54145 33885 54179
rect 33919 54176 33931 54179
rect 34054 54176 34060 54188
rect 33919 54148 34060 54176
rect 33919 54145 33931 54148
rect 33873 54139 33931 54145
rect 34054 54136 34060 54148
rect 34112 54136 34118 54188
rect 35161 54179 35219 54185
rect 35161 54145 35173 54179
rect 35207 54176 35219 54179
rect 35342 54176 35348 54188
rect 35207 54148 35348 54176
rect 35207 54145 35219 54148
rect 35161 54139 35219 54145
rect 35342 54136 35348 54148
rect 35400 54136 35406 54188
rect 39209 54179 39267 54185
rect 39209 54145 39221 54179
rect 39255 54145 39267 54179
rect 39209 54139 39267 54145
rect 30098 54108 30104 54120
rect 29748 54080 30104 54108
rect 30098 54068 30104 54080
rect 30156 54108 30162 54120
rect 30469 54111 30527 54117
rect 30469 54108 30481 54111
rect 30156 54080 30481 54108
rect 30156 54068 30162 54080
rect 30469 54077 30481 54080
rect 30515 54077 30527 54111
rect 30469 54071 30527 54077
rect 30745 54111 30803 54117
rect 30745 54077 30757 54111
rect 30791 54108 30803 54111
rect 31018 54108 31024 54120
rect 30791 54080 31024 54108
rect 30791 54077 30803 54080
rect 30745 54071 30803 54077
rect 30484 54040 30512 54071
rect 31018 54068 31024 54080
rect 31076 54068 31082 54120
rect 32214 54068 32220 54120
rect 32272 54108 32278 54120
rect 32401 54111 32459 54117
rect 32401 54108 32413 54111
rect 32272 54080 32413 54108
rect 32272 54068 32278 54080
rect 32401 54077 32413 54080
rect 32447 54077 32459 54111
rect 32401 54071 32459 54077
rect 32582 54068 32588 54120
rect 32640 54108 32646 54120
rect 33965 54111 34023 54117
rect 33965 54108 33977 54111
rect 32640 54080 33977 54108
rect 32640 54068 32646 54080
rect 33965 54077 33977 54080
rect 34011 54108 34023 54111
rect 34146 54108 34152 54120
rect 34011 54080 34152 54108
rect 34011 54077 34023 54080
rect 33965 54071 34023 54077
rect 34146 54068 34152 54080
rect 34204 54108 34210 54120
rect 34698 54108 34704 54120
rect 34204 54080 34704 54108
rect 34204 54068 34210 54080
rect 34698 54068 34704 54080
rect 34756 54068 34762 54120
rect 34790 54068 34796 54120
rect 34848 54108 34854 54120
rect 35069 54111 35127 54117
rect 35069 54108 35081 54111
rect 34848 54080 35081 54108
rect 34848 54068 34854 54080
rect 35069 54077 35081 54080
rect 35115 54077 35127 54111
rect 39224 54108 39252 54139
rect 39574 54136 39580 54188
rect 39632 54176 39638 54188
rect 39669 54179 39727 54185
rect 39669 54176 39681 54179
rect 39632 54148 39681 54176
rect 39632 54136 39638 54148
rect 39669 54145 39681 54148
rect 39715 54145 39727 54179
rect 40310 54176 40316 54188
rect 40271 54148 40316 54176
rect 39669 54139 39727 54145
rect 40310 54136 40316 54148
rect 40368 54136 40374 54188
rect 41138 54176 41144 54188
rect 41099 54148 41144 54176
rect 41138 54136 41144 54148
rect 41196 54136 41202 54188
rect 42610 54176 42616 54188
rect 42571 54148 42616 54176
rect 42610 54136 42616 54148
rect 42668 54136 42674 54188
rect 42889 54179 42947 54185
rect 42889 54145 42901 54179
rect 42935 54176 42947 54179
rect 42978 54176 42984 54188
rect 42935 54148 42984 54176
rect 42935 54145 42947 54148
rect 42889 54139 42947 54145
rect 42978 54136 42984 54148
rect 43036 54136 43042 54188
rect 43254 54136 43260 54188
rect 43312 54176 43318 54188
rect 43809 54179 43867 54185
rect 43809 54176 43821 54179
rect 43312 54148 43821 54176
rect 43312 54136 43318 54148
rect 43809 54145 43821 54148
rect 43855 54145 43867 54179
rect 43990 54176 43996 54188
rect 43951 54148 43996 54176
rect 43809 54139 43867 54145
rect 43990 54136 43996 54148
rect 44048 54136 44054 54188
rect 39942 54108 39948 54120
rect 39224 54080 39948 54108
rect 35069 54071 35127 54077
rect 39942 54068 39948 54080
rect 40000 54068 40006 54120
rect 41230 54108 41236 54120
rect 41191 54080 41236 54108
rect 41230 54068 41236 54080
rect 41288 54068 41294 54120
rect 43070 54068 43076 54120
rect 43128 54108 43134 54120
rect 43717 54111 43775 54117
rect 43717 54108 43729 54111
rect 43128 54080 43729 54108
rect 43128 54068 43134 54080
rect 43717 54077 43729 54080
rect 43763 54077 43775 54111
rect 43717 54071 43775 54077
rect 30484 54012 34928 54040
rect 33318 53932 33324 53984
rect 33376 53972 33382 53984
rect 34900 53981 34928 54012
rect 33689 53975 33747 53981
rect 33689 53972 33701 53975
rect 33376 53944 33701 53972
rect 33376 53932 33382 53944
rect 33689 53941 33701 53944
rect 33735 53941 33747 53975
rect 33689 53935 33747 53941
rect 34885 53975 34943 53981
rect 34885 53941 34897 53975
rect 34931 53941 34943 53975
rect 34885 53935 34943 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 27706 53728 27712 53780
rect 27764 53768 27770 53780
rect 27893 53771 27951 53777
rect 27893 53768 27905 53771
rect 27764 53740 27905 53768
rect 27764 53728 27770 53740
rect 27893 53737 27905 53740
rect 27939 53737 27951 53771
rect 27893 53731 27951 53737
rect 29730 53728 29736 53780
rect 29788 53768 29794 53780
rect 29917 53771 29975 53777
rect 29917 53768 29929 53771
rect 29788 53740 29929 53768
rect 29788 53728 29794 53740
rect 29917 53737 29929 53740
rect 29963 53737 29975 53771
rect 30742 53768 30748 53780
rect 30703 53740 30748 53768
rect 29917 53731 29975 53737
rect 30742 53728 30748 53740
rect 30800 53728 30806 53780
rect 31110 53728 31116 53780
rect 31168 53768 31174 53780
rect 31941 53771 31999 53777
rect 31941 53768 31953 53771
rect 31168 53740 31953 53768
rect 31168 53728 31174 53740
rect 31941 53737 31953 53740
rect 31987 53737 31999 53771
rect 31941 53731 31999 53737
rect 32861 53771 32919 53777
rect 32861 53737 32873 53771
rect 32907 53768 32919 53771
rect 33134 53768 33140 53780
rect 32907 53740 33140 53768
rect 32907 53737 32919 53740
rect 32861 53731 32919 53737
rect 26973 53703 27031 53709
rect 26973 53669 26985 53703
rect 27019 53700 27031 53703
rect 29181 53703 29239 53709
rect 29181 53700 29193 53703
rect 27019 53672 29193 53700
rect 27019 53669 27031 53672
rect 26973 53663 27031 53669
rect 29181 53669 29193 53672
rect 29227 53700 29239 53703
rect 30760 53700 30788 53728
rect 31389 53703 31447 53709
rect 31389 53700 31401 53703
rect 29227 53672 31401 53700
rect 29227 53669 29239 53672
rect 29181 53663 29239 53669
rect 31389 53669 31401 53672
rect 31435 53700 31447 53703
rect 31478 53700 31484 53712
rect 31435 53672 31484 53700
rect 31435 53669 31447 53672
rect 31389 53663 31447 53669
rect 31478 53660 31484 53672
rect 31536 53660 31542 53712
rect 30282 53632 30288 53644
rect 30243 53604 30288 53632
rect 30282 53592 30288 53604
rect 30340 53592 30346 53644
rect 30098 53564 30104 53576
rect 30059 53536 30104 53564
rect 30098 53524 30104 53536
rect 30156 53524 30162 53576
rect 32122 53564 32128 53576
rect 32083 53536 32128 53564
rect 32122 53524 32128 53536
rect 32180 53524 32186 53576
rect 32214 53524 32220 53576
rect 32272 53564 32278 53576
rect 32401 53567 32459 53573
rect 32401 53564 32413 53567
rect 32272 53536 32413 53564
rect 32272 53524 32278 53536
rect 32401 53533 32413 53536
rect 32447 53533 32459 53567
rect 32401 53527 32459 53533
rect 32309 53499 32367 53505
rect 32309 53465 32321 53499
rect 32355 53496 32367 53499
rect 32876 53496 32904 53731
rect 33134 53728 33140 53740
rect 33192 53728 33198 53780
rect 33778 53728 33784 53780
rect 33836 53768 33842 53780
rect 33873 53771 33931 53777
rect 33873 53768 33885 53771
rect 33836 53740 33885 53768
rect 33836 53728 33842 53740
rect 33873 53737 33885 53740
rect 33919 53737 33931 53771
rect 33873 53731 33931 53737
rect 34790 53728 34796 53780
rect 34848 53768 34854 53780
rect 34885 53771 34943 53777
rect 34885 53768 34897 53771
rect 34848 53740 34897 53768
rect 34848 53728 34854 53740
rect 34885 53737 34897 53740
rect 34931 53737 34943 53771
rect 34885 53731 34943 53737
rect 35253 53771 35311 53777
rect 35253 53737 35265 53771
rect 35299 53768 35311 53771
rect 35526 53768 35532 53780
rect 35299 53740 35532 53768
rect 35299 53737 35311 53740
rect 35253 53731 35311 53737
rect 35526 53728 35532 53740
rect 35584 53728 35590 53780
rect 35894 53768 35900 53780
rect 35855 53740 35900 53768
rect 35894 53728 35900 53740
rect 35952 53728 35958 53780
rect 40221 53771 40279 53777
rect 40221 53737 40233 53771
rect 40267 53768 40279 53771
rect 40310 53768 40316 53780
rect 40267 53740 40316 53768
rect 40267 53737 40279 53740
rect 40221 53731 40279 53737
rect 40310 53728 40316 53740
rect 40368 53728 40374 53780
rect 42058 53768 42064 53780
rect 42019 53740 42064 53768
rect 42058 53728 42064 53740
rect 42116 53728 42122 53780
rect 42245 53771 42303 53777
rect 42245 53737 42257 53771
rect 42291 53768 42303 53771
rect 42702 53768 42708 53780
rect 42291 53740 42708 53768
rect 42291 53737 42303 53740
rect 42245 53731 42303 53737
rect 42702 53728 42708 53740
rect 42760 53728 42766 53780
rect 39393 53703 39451 53709
rect 39393 53669 39405 53703
rect 39439 53700 39451 53703
rect 39942 53700 39948 53712
rect 39439 53672 39948 53700
rect 39439 53669 39451 53672
rect 39393 53663 39451 53669
rect 39942 53660 39948 53672
rect 40000 53700 40006 53712
rect 40773 53703 40831 53709
rect 40773 53700 40785 53703
rect 40000 53672 40785 53700
rect 40000 53660 40006 53672
rect 40773 53669 40785 53672
rect 40819 53700 40831 53703
rect 41325 53703 41383 53709
rect 41325 53700 41337 53703
rect 40819 53672 41337 53700
rect 40819 53669 40831 53672
rect 40773 53663 40831 53669
rect 41325 53669 41337 53672
rect 41371 53700 41383 53703
rect 41966 53700 41972 53712
rect 41371 53672 41972 53700
rect 41371 53669 41383 53672
rect 41325 53663 41383 53669
rect 41966 53660 41972 53672
rect 42024 53660 42030 53712
rect 33962 53632 33968 53644
rect 33060 53604 33968 53632
rect 33060 53573 33088 53604
rect 33962 53592 33968 53604
rect 34020 53592 34026 53644
rect 34698 53592 34704 53644
rect 34756 53632 34762 53644
rect 35345 53635 35403 53641
rect 35345 53632 35357 53635
rect 34756 53604 35357 53632
rect 34756 53592 34762 53604
rect 35345 53601 35357 53604
rect 35391 53601 35403 53635
rect 35345 53595 35403 53601
rect 33045 53567 33103 53573
rect 33045 53533 33057 53567
rect 33091 53533 33103 53567
rect 33318 53564 33324 53576
rect 33279 53536 33324 53564
rect 33045 53527 33103 53533
rect 33318 53524 33324 53536
rect 33376 53524 33382 53576
rect 34054 53564 34060 53576
rect 34015 53536 34060 53564
rect 34054 53524 34060 53536
rect 34112 53524 34118 53576
rect 34146 53524 34152 53576
rect 34204 53573 34210 53576
rect 34330 53573 34336 53576
rect 34204 53567 34217 53573
rect 34205 53564 34217 53567
rect 34277 53567 34336 53573
rect 34205 53536 34249 53564
rect 34205 53533 34217 53536
rect 34204 53527 34217 53533
rect 34277 53533 34289 53567
rect 34323 53533 34336 53567
rect 34277 53527 34336 53533
rect 34204 53524 34210 53527
rect 34330 53524 34336 53527
rect 34388 53524 34394 53576
rect 35069 53567 35127 53573
rect 35069 53533 35081 53567
rect 35115 53533 35127 53567
rect 35069 53527 35127 53533
rect 32355 53468 32904 53496
rect 33229 53499 33287 53505
rect 32355 53465 32367 53468
rect 32309 53459 32367 53465
rect 33229 53465 33241 53499
rect 33275 53496 33287 53499
rect 33778 53496 33784 53508
rect 33275 53468 33784 53496
rect 33275 53465 33287 53468
rect 33229 53459 33287 53465
rect 33778 53456 33784 53468
rect 33836 53456 33842 53508
rect 34072 53496 34100 53524
rect 35084 53496 35112 53527
rect 34072 53468 35112 53496
rect 42429 53499 42487 53505
rect 42429 53465 42441 53499
rect 42475 53496 42487 53499
rect 42978 53496 42984 53508
rect 42475 53468 42984 53496
rect 42475 53465 42487 53468
rect 42429 53459 42487 53465
rect 42978 53456 42984 53468
rect 43036 53456 43042 53508
rect 42229 53431 42287 53437
rect 42229 53397 42241 53431
rect 42275 53428 42287 53431
rect 42610 53428 42616 53440
rect 42275 53400 42616 53428
rect 42275 53397 42287 53400
rect 42229 53391 42287 53397
rect 42610 53388 42616 53400
rect 42668 53388 42674 53440
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 30466 53224 30472 53236
rect 30427 53196 30472 53224
rect 30466 53184 30472 53196
rect 30524 53184 30530 53236
rect 31478 53224 31484 53236
rect 31439 53196 31484 53224
rect 31478 53184 31484 53196
rect 31536 53184 31542 53236
rect 32398 53184 32404 53236
rect 32456 53224 32462 53236
rect 32769 53227 32827 53233
rect 32769 53224 32781 53227
rect 32456 53196 32781 53224
rect 32456 53184 32462 53196
rect 32769 53193 32781 53196
rect 32815 53224 32827 53227
rect 33321 53227 33379 53233
rect 33321 53224 33333 53227
rect 32815 53196 33333 53224
rect 32815 53193 32827 53196
rect 32769 53187 32827 53193
rect 33321 53193 33333 53196
rect 33367 53224 33379 53227
rect 33873 53227 33931 53233
rect 33873 53224 33885 53227
rect 33367 53196 33885 53224
rect 33367 53193 33379 53196
rect 33321 53187 33379 53193
rect 33873 53193 33885 53196
rect 33919 53224 33931 53227
rect 34425 53227 34483 53233
rect 34425 53224 34437 53227
rect 33919 53196 34437 53224
rect 33919 53193 33931 53196
rect 33873 53187 33931 53193
rect 34425 53193 34437 53196
rect 34471 53193 34483 53227
rect 39850 53224 39856 53236
rect 39811 53196 39856 53224
rect 34425 53187 34483 53193
rect 39850 53184 39856 53196
rect 39908 53184 39914 53236
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 32030 52640 32036 52692
rect 32088 52680 32094 52692
rect 32125 52683 32183 52689
rect 32125 52680 32137 52683
rect 32088 52652 32137 52680
rect 32088 52640 32094 52652
rect 32125 52649 32137 52652
rect 32171 52649 32183 52683
rect 32125 52643 32183 52649
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 34333 52071 34391 52077
rect 34333 52037 34345 52071
rect 34379 52068 34391 52071
rect 35986 52068 35992 52080
rect 34379 52040 35992 52068
rect 34379 52037 34391 52040
rect 34333 52031 34391 52037
rect 35986 52028 35992 52040
rect 36044 52028 36050 52080
rect 34146 51932 34152 51944
rect 34107 51904 34152 51932
rect 34146 51892 34152 51904
rect 34204 51892 34210 51944
rect 35710 51932 35716 51944
rect 35671 51904 35716 51932
rect 35710 51892 35716 51904
rect 35768 51892 35774 51944
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 34146 51592 34152 51604
rect 34107 51564 34152 51592
rect 34146 51552 34152 51564
rect 34204 51552 34210 51604
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 28994 8616 29000 8628
rect 26568 8588 29000 8616
rect 26568 8576 26574 8588
rect 28994 8576 29000 8588
rect 29052 8616 29058 8628
rect 29549 8619 29607 8625
rect 29549 8616 29561 8619
rect 29052 8588 29561 8616
rect 29052 8576 29058 8588
rect 29549 8585 29561 8588
rect 29595 8616 29607 8619
rect 29822 8616 29828 8628
rect 29595 8588 29828 8616
rect 29595 8585 29607 8588
rect 29549 8579 29607 8585
rect 29822 8576 29828 8588
rect 29880 8576 29886 8628
rect 30469 8483 30527 8489
rect 30469 8449 30481 8483
rect 30515 8449 30527 8483
rect 30469 8443 30527 8449
rect 30098 8236 30104 8288
rect 30156 8276 30162 8288
rect 30484 8276 30512 8443
rect 30561 8347 30619 8353
rect 30561 8313 30573 8347
rect 30607 8344 30619 8347
rect 30650 8344 30656 8356
rect 30607 8316 30656 8344
rect 30607 8313 30619 8316
rect 30561 8307 30619 8313
rect 30650 8304 30656 8316
rect 30708 8304 30714 8356
rect 30156 8248 30512 8276
rect 30156 8236 30162 8248
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 27522 7828 27528 7880
rect 27580 7868 27586 7880
rect 27801 7871 27859 7877
rect 27801 7868 27813 7871
rect 27580 7840 27813 7868
rect 27580 7828 27586 7840
rect 27801 7837 27813 7840
rect 27847 7837 27859 7871
rect 27801 7831 27859 7837
rect 28997 7871 29055 7877
rect 28997 7837 29009 7871
rect 29043 7868 29055 7871
rect 29917 7871 29975 7877
rect 29917 7868 29929 7871
rect 29043 7840 29929 7868
rect 29043 7837 29055 7840
rect 28997 7831 29055 7837
rect 29917 7837 29929 7840
rect 29963 7868 29975 7871
rect 30098 7868 30104 7880
rect 29963 7840 30104 7868
rect 29963 7837 29975 7840
rect 29917 7831 29975 7837
rect 30098 7828 30104 7840
rect 30156 7828 30162 7880
rect 30466 7868 30472 7880
rect 30427 7840 30472 7868
rect 30466 7828 30472 7840
rect 30524 7828 30530 7880
rect 31297 7871 31355 7877
rect 31297 7837 31309 7871
rect 31343 7837 31355 7871
rect 31297 7831 31355 7837
rect 30116 7800 30144 7828
rect 31312 7800 31340 7831
rect 30116 7772 31340 7800
rect 27614 7692 27620 7744
rect 27672 7732 27678 7744
rect 27893 7735 27951 7741
rect 27893 7732 27905 7735
rect 27672 7704 27905 7732
rect 27672 7692 27678 7704
rect 27893 7701 27905 7704
rect 27939 7701 27951 7735
rect 27893 7695 27951 7701
rect 29089 7735 29147 7741
rect 29089 7701 29101 7735
rect 29135 7732 29147 7735
rect 29362 7732 29368 7744
rect 29135 7704 29368 7732
rect 29135 7701 29147 7704
rect 29089 7695 29147 7701
rect 29362 7692 29368 7704
rect 29420 7692 29426 7744
rect 29546 7692 29552 7744
rect 29604 7732 29610 7744
rect 29825 7735 29883 7741
rect 29825 7732 29837 7735
rect 29604 7704 29837 7732
rect 29604 7692 29610 7704
rect 29825 7701 29837 7704
rect 29871 7701 29883 7735
rect 29825 7695 29883 7701
rect 31110 7692 31116 7744
rect 31168 7732 31174 7744
rect 31205 7735 31263 7741
rect 31205 7732 31217 7735
rect 31168 7704 31217 7732
rect 31168 7692 31174 7704
rect 31205 7701 31217 7704
rect 31251 7701 31263 7735
rect 31205 7695 31263 7701
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 29546 7460 29552 7472
rect 29507 7432 29552 7460
rect 29546 7420 29552 7432
rect 29604 7420 29610 7472
rect 28905 7327 28963 7333
rect 28905 7293 28917 7327
rect 28951 7324 28963 7327
rect 29365 7327 29423 7333
rect 29365 7324 29377 7327
rect 28951 7296 29377 7324
rect 28951 7293 28963 7296
rect 28905 7287 28963 7293
rect 29365 7293 29377 7296
rect 29411 7293 29423 7327
rect 30742 7324 30748 7336
rect 30703 7296 30748 7324
rect 29365 7287 29423 7293
rect 30742 7284 30748 7296
rect 30800 7284 30806 7336
rect 27338 7188 27344 7200
rect 27299 7160 27344 7188
rect 27338 7148 27344 7160
rect 27396 7148 27402 7200
rect 27982 7188 27988 7200
rect 27943 7160 27988 7188
rect 27982 7148 27988 7160
rect 28040 7148 28046 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 27338 6848 27344 6860
rect 27299 6820 27344 6848
rect 27338 6808 27344 6820
rect 27396 6808 27402 6860
rect 27525 6851 27583 6857
rect 27525 6817 27537 6851
rect 27571 6848 27583 6851
rect 27614 6848 27620 6860
rect 27571 6820 27620 6848
rect 27571 6817 27583 6820
rect 27525 6811 27583 6817
rect 27614 6808 27620 6820
rect 27672 6808 27678 6860
rect 28074 6848 28080 6860
rect 28035 6820 28080 6848
rect 28074 6808 28080 6820
rect 28132 6808 28138 6860
rect 31110 6848 31116 6860
rect 31071 6820 31116 6848
rect 31110 6808 31116 6820
rect 31168 6808 31174 6860
rect 31662 6848 31668 6860
rect 31623 6820 31668 6848
rect 31662 6808 31668 6820
rect 31720 6808 31726 6860
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6780 24915 6783
rect 25501 6783 25559 6789
rect 25501 6780 25513 6783
rect 24903 6752 25513 6780
rect 24903 6749 24915 6752
rect 24857 6743 24915 6749
rect 25501 6749 25513 6752
rect 25547 6780 25559 6783
rect 25547 6752 26280 6780
rect 25547 6749 25559 6752
rect 25501 6743 25559 6749
rect 25222 6604 25228 6656
rect 25280 6644 25286 6656
rect 26252 6653 26280 6752
rect 26418 6740 26424 6792
rect 26476 6780 26482 6792
rect 26697 6783 26755 6789
rect 26697 6780 26709 6783
rect 26476 6752 26709 6780
rect 26476 6740 26482 6752
rect 26697 6749 26709 6752
rect 26743 6749 26755 6783
rect 26697 6743 26755 6749
rect 29733 6783 29791 6789
rect 29733 6749 29745 6783
rect 29779 6780 29791 6783
rect 29822 6780 29828 6792
rect 29779 6752 29828 6780
rect 29779 6749 29791 6752
rect 29733 6743 29791 6749
rect 29822 6740 29828 6752
rect 29880 6740 29886 6792
rect 30926 6780 30932 6792
rect 30887 6752 30932 6780
rect 30926 6740 30932 6752
rect 30984 6740 30990 6792
rect 33781 6783 33839 6789
rect 33781 6749 33793 6783
rect 33827 6780 33839 6783
rect 35342 6780 35348 6792
rect 33827 6752 35348 6780
rect 33827 6749 33839 6752
rect 33781 6743 33839 6749
rect 35342 6740 35348 6752
rect 35400 6740 35406 6792
rect 30009 6715 30067 6721
rect 30009 6681 30021 6715
rect 30055 6712 30067 6715
rect 30098 6712 30104 6724
rect 30055 6684 30104 6712
rect 30055 6681 30067 6684
rect 30009 6675 30067 6681
rect 30098 6672 30104 6684
rect 30156 6672 30162 6724
rect 25409 6647 25467 6653
rect 25409 6644 25421 6647
rect 25280 6616 25421 6644
rect 25280 6604 25286 6616
rect 25409 6613 25421 6616
rect 25455 6613 25467 6647
rect 25409 6607 25467 6613
rect 26237 6647 26295 6653
rect 26237 6613 26249 6647
rect 26283 6644 26295 6647
rect 26510 6644 26516 6656
rect 26283 6616 26516 6644
rect 26283 6613 26295 6616
rect 26237 6607 26295 6613
rect 26510 6604 26516 6616
rect 26568 6604 26574 6656
rect 26789 6647 26847 6653
rect 26789 6613 26801 6647
rect 26835 6644 26847 6647
rect 27338 6644 27344 6656
rect 26835 6616 27344 6644
rect 26835 6613 26847 6616
rect 26789 6607 26847 6613
rect 27338 6604 27344 6616
rect 27396 6604 27402 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 29822 6400 29828 6452
rect 29880 6440 29886 6452
rect 32766 6440 32772 6452
rect 29880 6412 32772 6440
rect 29880 6400 29886 6412
rect 32766 6400 32772 6412
rect 32824 6440 32830 6452
rect 32953 6443 33011 6449
rect 32953 6440 32965 6443
rect 32824 6412 32965 6440
rect 32824 6400 32830 6412
rect 32953 6409 32965 6412
rect 32999 6409 33011 6443
rect 32953 6403 33011 6409
rect 29362 6372 29368 6384
rect 29323 6344 29368 6372
rect 29362 6332 29368 6344
rect 29420 6332 29426 6384
rect 26418 6304 26424 6316
rect 26379 6276 26424 6304
rect 26418 6264 26424 6276
rect 26476 6264 26482 6316
rect 26510 6264 26516 6316
rect 26568 6304 26574 6316
rect 27249 6307 27307 6313
rect 27249 6304 27261 6307
rect 26568 6276 27261 6304
rect 26568 6264 26574 6276
rect 27249 6273 27261 6276
rect 27295 6304 27307 6307
rect 28994 6304 29000 6316
rect 27295 6276 29000 6304
rect 27295 6273 27307 6276
rect 27249 6267 27307 6273
rect 28994 6264 29000 6276
rect 29052 6264 29058 6316
rect 30926 6264 30932 6316
rect 30984 6304 30990 6316
rect 31481 6307 31539 6313
rect 31481 6304 31493 6307
rect 30984 6276 31493 6304
rect 30984 6264 30990 6276
rect 31481 6273 31493 6276
rect 31527 6273 31539 6307
rect 31481 6267 31539 6273
rect 35342 6264 35348 6316
rect 35400 6304 35406 6316
rect 35400 6276 35445 6304
rect 35400 6264 35406 6276
rect 26436 6236 26464 6264
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 26436 6208 27445 6236
rect 27433 6205 27445 6208
rect 27479 6236 27491 6239
rect 27522 6236 27528 6248
rect 27479 6208 27528 6236
rect 27479 6205 27491 6208
rect 27433 6199 27491 6205
rect 27522 6196 27528 6208
rect 27580 6196 27586 6248
rect 29178 6236 29184 6248
rect 29139 6208 29184 6236
rect 29178 6196 29184 6208
rect 29236 6196 29242 6248
rect 29730 6236 29736 6248
rect 29691 6208 29736 6236
rect 29730 6196 29736 6208
rect 29788 6196 29794 6248
rect 33870 6236 33876 6248
rect 33831 6208 33876 6236
rect 33870 6196 33876 6208
rect 33928 6196 33934 6248
rect 35161 6239 35219 6245
rect 35161 6205 35173 6239
rect 35207 6205 35219 6239
rect 35161 6199 35219 6205
rect 35176 6168 35204 6199
rect 35618 6168 35624 6180
rect 35176 6140 35624 6168
rect 35618 6128 35624 6140
rect 35676 6128 35682 6180
rect 25038 6060 25044 6112
rect 25096 6100 25102 6112
rect 25409 6103 25467 6109
rect 25409 6100 25421 6103
rect 25096 6072 25421 6100
rect 25096 6060 25102 6072
rect 25409 6069 25421 6072
rect 25455 6069 25467 6103
rect 25409 6063 25467 6069
rect 26513 6103 26571 6109
rect 26513 6069 26525 6103
rect 26559 6100 26571 6103
rect 27522 6100 27528 6112
rect 26559 6072 27528 6100
rect 26559 6069 26571 6072
rect 26513 6063 26571 6069
rect 27522 6060 27528 6072
rect 27580 6060 27586 6112
rect 28721 6103 28779 6109
rect 28721 6069 28733 6103
rect 28767 6100 28779 6103
rect 29454 6100 29460 6112
rect 28767 6072 29460 6100
rect 28767 6069 28779 6072
rect 28721 6063 28779 6069
rect 29454 6060 29460 6072
rect 29512 6060 29518 6112
rect 32493 6103 32551 6109
rect 32493 6069 32505 6103
rect 32539 6100 32551 6103
rect 34146 6100 34152 6112
rect 32539 6072 34152 6100
rect 32539 6069 32551 6072
rect 32493 6063 32551 6069
rect 34146 6060 34152 6072
rect 34204 6060 34210 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 35618 5896 35624 5908
rect 35579 5868 35624 5896
rect 35618 5856 35624 5868
rect 35676 5856 35682 5908
rect 27982 5828 27988 5840
rect 27356 5800 27988 5828
rect 25038 5760 25044 5772
rect 24999 5732 25044 5760
rect 25038 5720 25044 5732
rect 25096 5720 25102 5772
rect 25222 5760 25228 5772
rect 25183 5732 25228 5760
rect 25222 5720 25228 5732
rect 25280 5720 25286 5772
rect 25958 5760 25964 5772
rect 25919 5732 25964 5760
rect 25958 5720 25964 5732
rect 26016 5720 26022 5772
rect 27356 5769 27384 5800
rect 27982 5788 27988 5800
rect 28040 5788 28046 5840
rect 27341 5763 27399 5769
rect 27341 5729 27353 5763
rect 27387 5729 27399 5763
rect 27522 5760 27528 5772
rect 27483 5732 27528 5760
rect 27341 5723 27399 5729
rect 27522 5720 27528 5732
rect 27580 5720 27586 5772
rect 27798 5760 27804 5772
rect 27759 5732 27804 5760
rect 27798 5720 27804 5732
rect 27856 5720 27862 5772
rect 30466 5760 30472 5772
rect 30427 5732 30472 5760
rect 30466 5720 30472 5732
rect 30524 5720 30530 5772
rect 30650 5760 30656 5772
rect 30611 5732 30656 5760
rect 30650 5720 30656 5732
rect 30708 5720 30714 5772
rect 31386 5760 31392 5772
rect 31347 5732 31392 5760
rect 31386 5720 31392 5732
rect 31444 5720 31450 5772
rect 35342 5760 35348 5772
rect 33704 5732 35348 5760
rect 29914 5652 29920 5704
rect 29972 5692 29978 5704
rect 30009 5695 30067 5701
rect 30009 5692 30021 5695
rect 29972 5664 30021 5692
rect 29972 5652 29978 5664
rect 30009 5661 30021 5664
rect 30055 5661 30067 5695
rect 32766 5692 32772 5704
rect 32727 5664 32772 5692
rect 30009 5655 30067 5661
rect 32766 5652 32772 5664
rect 32824 5652 32830 5704
rect 33704 5701 33732 5732
rect 35342 5720 35348 5732
rect 35400 5760 35406 5772
rect 35400 5732 35756 5760
rect 35400 5720 35406 5732
rect 33045 5695 33103 5701
rect 33045 5661 33057 5695
rect 33091 5692 33103 5695
rect 33689 5695 33747 5701
rect 33689 5692 33701 5695
rect 33091 5664 33701 5692
rect 33091 5661 33103 5664
rect 33045 5655 33103 5661
rect 33689 5661 33701 5664
rect 33735 5661 33747 5695
rect 33689 5655 33747 5661
rect 34514 5652 34520 5704
rect 34572 5692 34578 5704
rect 35728 5701 35756 5732
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34572 5664 34897 5692
rect 34572 5652 34578 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5692 35771 5695
rect 36357 5695 36415 5701
rect 36357 5692 36369 5695
rect 35759 5664 36369 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 36357 5661 36369 5664
rect 36403 5661 36415 5695
rect 36357 5655 36415 5661
rect 33781 5559 33839 5565
rect 33781 5525 33793 5559
rect 33827 5556 33839 5559
rect 33962 5556 33968 5568
rect 33827 5528 33968 5556
rect 33827 5525 33839 5528
rect 33781 5519 33839 5525
rect 33962 5516 33968 5528
rect 34020 5516 34026 5568
rect 36262 5556 36268 5568
rect 36223 5528 36268 5556
rect 36262 5516 36268 5528
rect 36320 5516 36326 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 27338 5284 27344 5296
rect 27299 5256 27344 5284
rect 27338 5244 27344 5256
rect 27396 5244 27402 5296
rect 33962 5284 33968 5296
rect 33923 5256 33968 5284
rect 33962 5244 33968 5256
rect 34020 5244 34026 5296
rect 36262 5284 36268 5296
rect 36223 5256 36268 5284
rect 36262 5244 36268 5256
rect 36320 5244 36326 5296
rect 29454 5216 29460 5228
rect 29415 5188 29460 5216
rect 29454 5176 29460 5188
rect 29512 5176 29518 5228
rect 34146 5176 34152 5228
rect 34204 5216 34210 5228
rect 34204 5188 34249 5216
rect 34204 5176 34210 5188
rect 26605 5151 26663 5157
rect 26605 5117 26617 5151
rect 26651 5148 26663 5151
rect 27157 5151 27215 5157
rect 27157 5148 27169 5151
rect 26651 5120 27169 5148
rect 26651 5117 26663 5120
rect 26605 5111 26663 5117
rect 27157 5117 27169 5120
rect 27203 5117 27215 5151
rect 27706 5148 27712 5160
rect 27667 5120 27712 5148
rect 27157 5111 27215 5117
rect 27706 5108 27712 5120
rect 27764 5108 27770 5160
rect 29638 5148 29644 5160
rect 29599 5120 29644 5148
rect 29638 5108 29644 5120
rect 29696 5108 29702 5160
rect 30374 5148 30380 5160
rect 30335 5120 30380 5148
rect 30374 5108 30380 5120
rect 30432 5108 30438 5160
rect 32490 5148 32496 5160
rect 32451 5120 32496 5148
rect 32490 5108 32496 5120
rect 32548 5108 32554 5160
rect 34698 5148 34704 5160
rect 34659 5120 34704 5148
rect 34698 5108 34704 5120
rect 34756 5108 34762 5160
rect 36446 5148 36452 5160
rect 36407 5120 36452 5148
rect 36446 5108 36452 5120
rect 36504 5108 36510 5160
rect 23658 4972 23664 5024
rect 23716 5012 23722 5024
rect 23753 5015 23811 5021
rect 23753 5012 23765 5015
rect 23716 4984 23765 5012
rect 23716 4972 23722 4984
rect 23753 4981 23765 4984
rect 23799 4981 23811 5015
rect 24670 5012 24676 5024
rect 24631 4984 24676 5012
rect 23753 4975 23811 4981
rect 24670 4972 24676 4984
rect 24728 4972 24734 5024
rect 25314 5012 25320 5024
rect 25275 4984 25320 5012
rect 25314 4972 25320 4984
rect 25372 4972 25378 5024
rect 25961 5015 26019 5021
rect 25961 4981 25973 5015
rect 26007 5012 26019 5015
rect 27338 5012 27344 5024
rect 26007 4984 27344 5012
rect 26007 4981 26019 4984
rect 25961 4975 26019 4981
rect 27338 4972 27344 4984
rect 27396 4972 27402 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 26418 4808 26424 4820
rect 24688 4780 26424 4808
rect 23385 4743 23443 4749
rect 23385 4709 23397 4743
rect 23431 4740 23443 4743
rect 23842 4740 23848 4752
rect 23431 4712 23848 4740
rect 23431 4709 23443 4712
rect 23385 4703 23443 4709
rect 23842 4700 23848 4712
rect 23900 4700 23906 4752
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 21545 4607 21603 4613
rect 21545 4604 21557 4607
rect 21508 4576 21557 4604
rect 21508 4564 21514 4576
rect 21545 4573 21557 4576
rect 21591 4573 21603 4607
rect 21545 4567 21603 4573
rect 22278 4564 22284 4616
rect 22336 4604 22342 4616
rect 22373 4607 22431 4613
rect 22373 4604 22385 4607
rect 22336 4576 22385 4604
rect 22336 4564 22342 4576
rect 22373 4573 22385 4576
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 23474 4564 23480 4616
rect 23532 4604 23538 4616
rect 24688 4613 24716 4780
rect 26418 4768 26424 4780
rect 26476 4768 26482 4820
rect 29178 4808 29184 4820
rect 29139 4780 29184 4808
rect 29178 4768 29184 4780
rect 29236 4768 29242 4820
rect 36357 4811 36415 4817
rect 36357 4777 36369 4811
rect 36403 4808 36415 4811
rect 36446 4808 36452 4820
rect 36403 4780 36452 4808
rect 36403 4777 36415 4780
rect 36357 4771 36415 4777
rect 36446 4768 36452 4780
rect 36504 4768 36510 4820
rect 25501 4743 25559 4749
rect 25501 4709 25513 4743
rect 25547 4740 25559 4743
rect 26878 4740 26884 4752
rect 25547 4712 26884 4740
rect 25547 4709 25559 4712
rect 25501 4703 25559 4709
rect 26878 4700 26884 4712
rect 26936 4700 26942 4752
rect 25314 4632 25320 4684
rect 25372 4672 25378 4684
rect 26605 4675 26663 4681
rect 26605 4672 26617 4675
rect 25372 4644 26617 4672
rect 25372 4632 25378 4644
rect 26605 4641 26617 4644
rect 26651 4641 26663 4675
rect 27614 4672 27620 4684
rect 27575 4644 27620 4672
rect 26605 4635 26663 4641
rect 27614 4632 27620 4644
rect 27672 4632 27678 4684
rect 29914 4672 29920 4684
rect 29875 4644 29920 4672
rect 29914 4632 29920 4644
rect 29972 4632 29978 4684
rect 30558 4672 30564 4684
rect 30519 4644 30564 4672
rect 30558 4632 30564 4644
rect 30616 4632 30622 4684
rect 32674 4672 32680 4684
rect 32635 4644 32680 4672
rect 32674 4632 32680 4644
rect 32732 4632 32738 4684
rect 34057 4675 34115 4681
rect 34057 4641 34069 4675
rect 34103 4672 34115 4675
rect 34514 4672 34520 4684
rect 34103 4644 34520 4672
rect 34103 4641 34115 4644
rect 34057 4635 34115 4641
rect 34514 4632 34520 4644
rect 34572 4632 34578 4684
rect 23845 4607 23903 4613
rect 23845 4604 23857 4607
rect 23532 4576 23857 4604
rect 23532 4564 23538 4576
rect 23845 4573 23857 4576
rect 23891 4604 23903 4607
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 23891 4576 24685 4604
rect 23891 4573 23903 4576
rect 23845 4567 23903 4573
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 26142 4604 26148 4616
rect 26103 4576 26148 4604
rect 24673 4567 24731 4573
rect 26142 4564 26148 4576
rect 26200 4564 26206 4616
rect 35069 4607 35127 4613
rect 35069 4573 35081 4607
rect 35115 4604 35127 4607
rect 35342 4604 35348 4616
rect 35115 4576 35348 4604
rect 35115 4573 35127 4576
rect 35069 4567 35127 4573
rect 35342 4564 35348 4576
rect 35400 4564 35406 4616
rect 35526 4604 35532 4616
rect 35487 4576 35532 4604
rect 35526 4564 35532 4576
rect 35584 4564 35590 4616
rect 36814 4604 36820 4616
rect 36775 4576 36820 4604
rect 36814 4564 36820 4576
rect 36872 4564 36878 4616
rect 23937 4539 23995 4545
rect 23937 4505 23949 4539
rect 23983 4536 23995 4539
rect 26789 4539 26847 4545
rect 26789 4536 26801 4539
rect 23983 4508 26801 4536
rect 23983 4505 23995 4508
rect 23937 4499 23995 4505
rect 26789 4505 26801 4508
rect 26835 4505 26847 4539
rect 26789 4499 26847 4505
rect 30101 4539 30159 4545
rect 30101 4505 30113 4539
rect 30147 4536 30159 4539
rect 30466 4536 30472 4548
rect 30147 4508 30472 4536
rect 30147 4505 30159 4508
rect 30101 4499 30159 4505
rect 30466 4496 30472 4508
rect 30524 4496 30530 4548
rect 33873 4539 33931 4545
rect 33873 4505 33885 4539
rect 33919 4536 33931 4539
rect 34977 4539 35035 4545
rect 34977 4536 34989 4539
rect 33919 4508 34989 4536
rect 33919 4505 33931 4508
rect 33873 4499 33931 4505
rect 34977 4505 34989 4508
rect 35023 4505 35035 4539
rect 34977 4499 35035 4505
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4468 24823 4471
rect 26050 4468 26056 4480
rect 24811 4440 26056 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 26050 4428 26056 4440
rect 26108 4428 26114 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 26142 4224 26148 4276
rect 26200 4264 26206 4276
rect 26200 4236 29960 4264
rect 26200 4224 26206 4236
rect 23474 4128 23480 4140
rect 23435 4100 23480 4128
rect 23474 4088 23480 4100
rect 23532 4088 23538 4140
rect 24670 4088 24676 4140
rect 24728 4128 24734 4140
rect 24765 4131 24823 4137
rect 24765 4128 24777 4131
rect 24728 4100 24777 4128
rect 24728 4088 24734 4100
rect 24765 4097 24777 4100
rect 24811 4097 24823 4131
rect 24765 4091 24823 4097
rect 26878 4088 26884 4140
rect 26936 4128 26942 4140
rect 29932 4137 29960 4236
rect 27617 4131 27675 4137
rect 27617 4128 27629 4131
rect 26936 4100 27629 4128
rect 26936 4088 26942 4100
rect 27617 4097 27629 4100
rect 27663 4097 27675 4131
rect 27617 4091 27675 4097
rect 29917 4131 29975 4137
rect 29917 4097 29929 4131
rect 29963 4097 29975 4131
rect 29917 4091 29975 4097
rect 34606 4088 34612 4140
rect 34664 4128 34670 4140
rect 34977 4131 35035 4137
rect 34977 4128 34989 4131
rect 34664 4100 34989 4128
rect 34664 4088 34670 4100
rect 34977 4097 34989 4100
rect 35023 4097 35035 4131
rect 34977 4091 35035 4097
rect 35342 4088 35348 4140
rect 35400 4128 35406 4140
rect 35618 4128 35624 4140
rect 35400 4100 35624 4128
rect 35400 4088 35406 4100
rect 35618 4088 35624 4100
rect 35676 4128 35682 4140
rect 35805 4131 35863 4137
rect 35805 4128 35817 4131
rect 35676 4100 35817 4128
rect 35676 4088 35682 4100
rect 35805 4097 35817 4100
rect 35851 4128 35863 4131
rect 37366 4128 37372 4140
rect 35851 4100 37372 4128
rect 35851 4097 35863 4100
rect 35805 4091 35863 4097
rect 37366 4088 37372 4100
rect 37424 4088 37430 4140
rect 23569 4063 23627 4069
rect 23569 4029 23581 4063
rect 23615 4060 23627 4063
rect 24949 4063 25007 4069
rect 24949 4060 24961 4063
rect 23615 4032 24961 4060
rect 23615 4029 23627 4032
rect 23569 4023 23627 4029
rect 24949 4029 24961 4032
rect 24995 4029 25007 4063
rect 26418 4060 26424 4072
rect 26379 4032 26424 4060
rect 24949 4023 25007 4029
rect 26418 4020 26424 4032
rect 26476 4020 26482 4072
rect 27801 4063 27859 4069
rect 27801 4029 27813 4063
rect 27847 4029 27859 4063
rect 28350 4060 28356 4072
rect 28311 4032 28356 4060
rect 27801 4023 27859 4029
rect 22373 3995 22431 4001
rect 22373 3961 22385 3995
rect 22419 3992 22431 3995
rect 23106 3992 23112 4004
rect 22419 3964 23112 3992
rect 22419 3961 22431 3964
rect 22373 3955 22431 3961
rect 23106 3952 23112 3964
rect 23164 3952 23170 4004
rect 25314 3992 25320 4004
rect 24228 3964 25320 3992
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17405 3927 17463 3933
rect 17405 3924 17417 3927
rect 17368 3896 17417 3924
rect 17368 3884 17374 3896
rect 17405 3893 17417 3896
rect 17451 3893 17463 3927
rect 17405 3887 17463 3893
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 19613 3927 19671 3933
rect 19613 3924 19625 3927
rect 19484 3896 19625 3924
rect 19484 3884 19490 3896
rect 19613 3893 19625 3896
rect 19659 3893 19671 3927
rect 19613 3887 19671 3893
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 20441 3927 20499 3933
rect 20441 3924 20453 3927
rect 20404 3896 20453 3924
rect 20404 3884 20410 3896
rect 20441 3893 20453 3896
rect 20487 3893 20499 3927
rect 20441 3887 20499 3893
rect 21453 3927 21511 3933
rect 21453 3893 21465 3927
rect 21499 3924 21511 3927
rect 22002 3924 22008 3936
rect 21499 3896 22008 3924
rect 21499 3893 21511 3896
rect 21453 3887 21511 3893
rect 22002 3884 22008 3896
rect 22060 3884 22066 3936
rect 23017 3927 23075 3933
rect 23017 3893 23029 3927
rect 23063 3924 23075 3927
rect 24228 3924 24256 3964
rect 25314 3952 25320 3964
rect 25372 3952 25378 4004
rect 26050 3952 26056 4004
rect 26108 3992 26114 4004
rect 27816 3992 27844 4023
rect 28350 4020 28356 4032
rect 28408 4020 28414 4072
rect 30101 4063 30159 4069
rect 30101 4029 30113 4063
rect 30147 4029 30159 4063
rect 30834 4060 30840 4072
rect 30795 4032 30840 4060
rect 30101 4023 30159 4029
rect 26108 3964 27844 3992
rect 26108 3952 26114 3964
rect 23063 3896 24256 3924
rect 24305 3927 24363 3933
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 24305 3893 24317 3927
rect 24351 3924 24363 3927
rect 25866 3924 25872 3936
rect 24351 3896 25872 3924
rect 24351 3893 24363 3896
rect 24305 3887 24363 3893
rect 25866 3884 25872 3896
rect 25924 3884 25930 3936
rect 30116 3924 30144 4023
rect 30834 4020 30840 4032
rect 30892 4020 30898 4072
rect 33042 4060 33048 4072
rect 33003 4032 33048 4060
rect 33042 4020 33048 4032
rect 33100 4020 33106 4072
rect 34333 4063 34391 4069
rect 34333 4029 34345 4063
rect 34379 4029 34391 4063
rect 34333 4023 34391 4029
rect 34517 4063 34575 4069
rect 34517 4029 34529 4063
rect 34563 4060 34575 4063
rect 35526 4060 35532 4072
rect 34563 4032 35532 4060
rect 34563 4029 34575 4032
rect 34517 4023 34575 4029
rect 34348 3992 34376 4023
rect 35526 4020 35532 4032
rect 35584 4020 35590 4072
rect 37461 4063 37519 4069
rect 37461 4060 37473 4063
rect 35820 4032 37473 4060
rect 35820 4004 35848 4032
rect 37461 4029 37473 4032
rect 37507 4029 37519 4063
rect 37461 4023 37519 4029
rect 35713 3995 35771 4001
rect 35713 3992 35725 3995
rect 34348 3964 35725 3992
rect 35713 3961 35725 3964
rect 35759 3961 35771 3995
rect 35713 3955 35771 3961
rect 35802 3952 35808 4004
rect 35860 3952 35866 4004
rect 37182 3952 37188 4004
rect 37240 3992 37246 4004
rect 38105 3995 38163 4001
rect 38105 3992 38117 3995
rect 37240 3964 38117 3992
rect 37240 3952 37246 3964
rect 38105 3961 38117 3964
rect 38151 3961 38163 3995
rect 38105 3955 38163 3961
rect 35069 3927 35127 3933
rect 35069 3924 35081 3927
rect 30116 3896 35081 3924
rect 35069 3893 35081 3896
rect 35115 3893 35127 3927
rect 35069 3887 35127 3893
rect 35434 3884 35440 3936
rect 35492 3924 35498 3936
rect 36265 3927 36323 3933
rect 36265 3924 36277 3927
rect 35492 3896 36277 3924
rect 35492 3884 35498 3896
rect 36265 3893 36277 3896
rect 36311 3893 36323 3927
rect 36265 3887 36323 3893
rect 38286 3884 38292 3936
rect 38344 3924 38350 3936
rect 38749 3927 38807 3933
rect 38749 3924 38761 3927
rect 38344 3896 38761 3924
rect 38344 3884 38350 3896
rect 38749 3893 38761 3896
rect 38795 3893 38807 3927
rect 38749 3887 38807 3893
rect 39390 3884 39396 3936
rect 39448 3924 39454 3936
rect 39485 3927 39543 3933
rect 39485 3924 39497 3927
rect 39448 3896 39497 3924
rect 39448 3884 39454 3896
rect 39485 3893 39497 3896
rect 39531 3893 39543 3927
rect 39485 3887 39543 3893
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 24486 3720 24492 3732
rect 22143 3692 24492 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 24486 3680 24492 3692
rect 24544 3680 24550 3732
rect 29638 3680 29644 3732
rect 29696 3720 29702 3732
rect 29825 3723 29883 3729
rect 29825 3720 29837 3723
rect 29696 3692 29837 3720
rect 29696 3680 29702 3692
rect 29825 3689 29837 3692
rect 29871 3689 29883 3723
rect 30466 3720 30472 3732
rect 30427 3692 30472 3720
rect 29825 3683 29883 3689
rect 30466 3680 30472 3692
rect 30524 3680 30530 3732
rect 34146 3680 34152 3732
rect 34204 3720 34210 3732
rect 34698 3720 34704 3732
rect 34204 3692 34704 3720
rect 34204 3680 34210 3692
rect 34698 3680 34704 3692
rect 34756 3680 34762 3732
rect 35526 3680 35532 3732
rect 35584 3720 35590 3732
rect 37829 3723 37887 3729
rect 37829 3720 37841 3723
rect 35584 3692 37841 3720
rect 35584 3680 35590 3692
rect 37829 3689 37841 3692
rect 37875 3689 37887 3723
rect 37829 3683 37887 3689
rect 21453 3655 21511 3661
rect 21453 3621 21465 3655
rect 21499 3652 21511 3655
rect 22830 3652 22836 3664
rect 21499 3624 22836 3652
rect 21499 3621 21511 3624
rect 21453 3615 21511 3621
rect 22830 3612 22836 3624
rect 22888 3612 22894 3664
rect 25682 3652 25688 3664
rect 23492 3624 25688 3652
rect 20809 3587 20867 3593
rect 20809 3553 20821 3587
rect 20855 3584 20867 3587
rect 21726 3584 21732 3596
rect 20855 3556 21732 3584
rect 20855 3553 20867 3556
rect 20809 3547 20867 3553
rect 21726 3544 21732 3556
rect 21784 3544 21790 3596
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3584 22799 3587
rect 23492 3584 23520 3624
rect 25682 3612 25688 3624
rect 25740 3612 25746 3664
rect 25774 3612 25780 3664
rect 25832 3652 25838 3664
rect 34606 3652 34612 3664
rect 25832 3624 29960 3652
rect 25832 3612 25838 3624
rect 22787 3556 23520 3584
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 23566 3544 23572 3596
rect 23624 3584 23630 3596
rect 25225 3587 25283 3593
rect 25225 3584 25237 3587
rect 23624 3556 25237 3584
rect 23624 3544 23630 3556
rect 25225 3553 25237 3556
rect 25271 3553 25283 3587
rect 26694 3584 26700 3596
rect 26655 3556 26700 3584
rect 25225 3547 25283 3553
rect 26694 3544 26700 3556
rect 26752 3544 26758 3596
rect 27338 3584 27344 3596
rect 27299 3556 27344 3584
rect 27338 3544 27344 3556
rect 27396 3544 27402 3596
rect 28902 3584 28908 3596
rect 28863 3556 28908 3584
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8996 3488 9137 3516
rect 8996 3476 9002 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10045 3519 10103 3525
rect 10045 3516 10057 3519
rect 10008 3488 10057 3516
rect 10008 3476 10014 3488
rect 10045 3485 10057 3488
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 10778 3476 10784 3528
rect 10836 3516 10842 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10836 3488 10885 3516
rect 10836 3476 10842 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 11606 3476 11612 3528
rect 11664 3516 11670 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11664 3488 11713 3516
rect 11664 3476 11670 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12492 3488 12541 3516
rect 12492 3476 12498 3488
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 13320 3488 13369 3516
rect 13320 3476 13326 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 14090 3476 14096 3528
rect 14148 3516 14154 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14148 3488 14289 3516
rect 14148 3476 14154 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14976 3488 15025 3516
rect 14976 3476 14982 3488
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 15746 3476 15752 3528
rect 15804 3516 15810 3528
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15804 3488 15853 3516
rect 15804 3476 15810 3488
rect 15841 3485 15853 3488
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16632 3488 16681 3516
rect 16632 3476 16638 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 17586 3516 17592 3528
rect 17547 3488 17592 3516
rect 16669 3479 16727 3485
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 18233 3519 18291 3525
rect 18233 3485 18245 3519
rect 18279 3516 18291 3519
rect 18414 3516 18420 3528
rect 18279 3488 18420 3516
rect 18279 3485 18291 3488
rect 18233 3479 18291 3485
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 19242 3516 19248 3528
rect 18923 3488 19248 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20622 3516 20628 3528
rect 20211 3488 20628 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 23400 3448 23428 3479
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23532 3488 23857 3516
rect 23532 3476 23538 3488
rect 23845 3485 23857 3488
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 23934 3476 23940 3528
rect 23992 3516 23998 3528
rect 29932 3525 29960 3624
rect 30576 3624 34612 3652
rect 25041 3519 25099 3525
rect 25041 3516 25053 3519
rect 23992 3488 25053 3516
rect 23992 3476 23998 3488
rect 25041 3485 25053 3488
rect 25087 3485 25099 3519
rect 25041 3479 25099 3485
rect 29917 3519 29975 3525
rect 29917 3485 29929 3519
rect 29963 3516 29975 3519
rect 30098 3516 30104 3528
rect 29963 3488 30104 3516
rect 29963 3485 29975 3488
rect 29917 3479 29975 3485
rect 30098 3476 30104 3488
rect 30156 3516 30162 3528
rect 30576 3525 30604 3624
rect 34606 3612 34612 3624
rect 34664 3612 34670 3664
rect 36906 3612 36912 3664
rect 36964 3652 36970 3664
rect 38473 3655 38531 3661
rect 38473 3652 38485 3655
rect 36964 3624 38485 3652
rect 36964 3612 36970 3624
rect 38473 3621 38485 3624
rect 38519 3621 38531 3655
rect 38473 3615 38531 3621
rect 39114 3612 39120 3664
rect 39172 3652 39178 3664
rect 40037 3655 40095 3661
rect 40037 3652 40049 3655
rect 39172 3624 40049 3652
rect 39172 3612 39178 3624
rect 40037 3621 40049 3624
rect 40083 3621 40095 3655
rect 40037 3615 40095 3621
rect 41046 3612 41052 3664
rect 41104 3652 41110 3664
rect 41969 3655 42027 3661
rect 41969 3652 41981 3655
rect 41104 3624 41981 3652
rect 41104 3612 41110 3624
rect 41969 3621 41981 3624
rect 42015 3621 42027 3655
rect 41969 3615 42027 3621
rect 45186 3612 45192 3664
rect 45244 3652 45250 3664
rect 45833 3655 45891 3661
rect 45833 3652 45845 3655
rect 45244 3624 45845 3652
rect 45244 3612 45250 3624
rect 45833 3621 45845 3624
rect 45879 3621 45891 3655
rect 45833 3615 45891 3621
rect 47118 3612 47124 3664
rect 47176 3652 47182 3664
rect 47765 3655 47823 3661
rect 47765 3652 47777 3655
rect 47176 3624 47777 3652
rect 47176 3612 47182 3624
rect 47765 3621 47777 3624
rect 47811 3621 47823 3655
rect 47765 3615 47823 3621
rect 36740 3596 36860 3600
rect 32214 3584 32220 3596
rect 32175 3556 32220 3584
rect 32214 3544 32220 3556
rect 32272 3544 32278 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 36740 3593 36820 3596
rect 34885 3587 34943 3593
rect 34885 3584 34897 3587
rect 33652 3556 34897 3584
rect 33652 3544 33658 3556
rect 34885 3553 34897 3556
rect 34931 3553 34943 3587
rect 34885 3547 34943 3553
rect 36725 3587 36820 3593
rect 36725 3553 36737 3587
rect 36771 3572 36820 3587
rect 36771 3553 36783 3572
rect 36725 3547 36783 3553
rect 36814 3544 36820 3572
rect 36872 3544 36878 3596
rect 39942 3544 39948 3596
rect 40000 3584 40006 3596
rect 40681 3587 40739 3593
rect 40681 3584 40693 3587
rect 40000 3556 40693 3584
rect 40000 3544 40006 3556
rect 40681 3553 40693 3556
rect 40727 3553 40739 3587
rect 40681 3547 40739 3553
rect 41874 3544 41880 3596
rect 41932 3584 41938 3596
rect 42613 3587 42671 3593
rect 42613 3584 42625 3587
rect 41932 3556 42625 3584
rect 41932 3544 41938 3556
rect 42613 3553 42625 3556
rect 42659 3553 42671 3587
rect 42613 3547 42671 3553
rect 42978 3544 42984 3596
rect 43036 3584 43042 3596
rect 43901 3587 43959 3593
rect 43901 3584 43913 3587
rect 43036 3556 43913 3584
rect 43036 3544 43042 3556
rect 43901 3553 43913 3556
rect 43947 3553 43959 3587
rect 43901 3547 43959 3553
rect 30561 3519 30619 3525
rect 30561 3516 30573 3519
rect 30156 3488 30573 3516
rect 30156 3476 30162 3488
rect 30561 3485 30573 3488
rect 30607 3485 30619 3519
rect 30561 3479 30619 3485
rect 33413 3519 33471 3525
rect 33413 3485 33425 3519
rect 33459 3516 33471 3519
rect 33873 3519 33931 3525
rect 33873 3516 33885 3519
rect 33459 3488 33885 3516
rect 33459 3485 33471 3488
rect 33413 3479 33471 3485
rect 33873 3485 33885 3488
rect 33919 3485 33931 3519
rect 37366 3516 37372 3528
rect 37327 3488 37372 3516
rect 33873 3479 33931 3485
rect 37366 3476 37372 3488
rect 37424 3476 37430 3528
rect 39117 3519 39175 3525
rect 39117 3485 39129 3519
rect 39163 3485 39175 3519
rect 39117 3479 39175 3485
rect 24762 3448 24768 3460
rect 23400 3420 24768 3448
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 27525 3451 27583 3457
rect 27525 3448 27537 3451
rect 26206 3420 27537 3448
rect 23937 3383 23995 3389
rect 23937 3349 23949 3383
rect 23983 3380 23995 3383
rect 26206 3380 26234 3420
rect 27525 3417 27537 3420
rect 27571 3417 27583 3451
rect 27525 3411 27583 3417
rect 30006 3408 30012 3460
rect 30064 3448 30070 3460
rect 30742 3448 30748 3460
rect 30064 3420 30748 3448
rect 30064 3408 30070 3420
rect 30742 3408 30748 3420
rect 30800 3408 30806 3460
rect 33229 3451 33287 3457
rect 33229 3417 33241 3451
rect 33275 3448 33287 3451
rect 34606 3448 34612 3460
rect 33275 3420 34612 3448
rect 33275 3417 33287 3420
rect 33229 3411 33287 3417
rect 34606 3408 34612 3420
rect 34664 3408 34670 3460
rect 36541 3451 36599 3457
rect 36541 3417 36553 3451
rect 36587 3448 36599 3451
rect 37277 3451 37335 3457
rect 37277 3448 37289 3451
rect 36587 3420 37289 3448
rect 36587 3417 36599 3420
rect 36541 3411 36599 3417
rect 37277 3417 37289 3420
rect 37323 3417 37335 3451
rect 37277 3411 37335 3417
rect 37642 3408 37648 3460
rect 37700 3448 37706 3460
rect 39132 3448 39160 3479
rect 40494 3476 40500 3528
rect 40552 3516 40558 3528
rect 41325 3519 41383 3525
rect 41325 3516 41337 3519
rect 40552 3488 41337 3516
rect 40552 3476 40558 3488
rect 41325 3485 41337 3488
rect 41371 3485 41383 3519
rect 41325 3479 41383 3485
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 43257 3519 43315 3525
rect 43257 3516 43269 3519
rect 42484 3488 43269 3516
rect 42484 3476 42490 3488
rect 43257 3485 43269 3488
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 44358 3476 44364 3528
rect 44416 3516 44422 3528
rect 45189 3519 45247 3525
rect 45189 3516 45201 3519
rect 44416 3488 45201 3516
rect 44416 3476 44422 3488
rect 45189 3485 45201 3488
rect 45235 3485 45247 3519
rect 45189 3479 45247 3485
rect 45738 3476 45744 3528
rect 45796 3516 45802 3528
rect 46477 3519 46535 3525
rect 46477 3516 46489 3519
rect 45796 3488 46489 3516
rect 45796 3476 45802 3488
rect 46477 3485 46489 3488
rect 46523 3485 46535 3519
rect 46477 3479 46535 3485
rect 47121 3519 47179 3525
rect 47121 3485 47133 3519
rect 47167 3485 47179 3519
rect 47121 3479 47179 3485
rect 37700 3420 39160 3448
rect 37700 3408 37706 3420
rect 46290 3408 46296 3460
rect 46348 3448 46354 3460
rect 47136 3448 47164 3479
rect 47946 3476 47952 3528
rect 48004 3516 48010 3528
rect 48409 3519 48467 3525
rect 48409 3516 48421 3519
rect 48004 3488 48421 3516
rect 48004 3476 48010 3488
rect 48409 3485 48421 3488
rect 48455 3485 48467 3519
rect 48409 3479 48467 3485
rect 49050 3476 49056 3528
rect 49108 3516 49114 3528
rect 49145 3519 49203 3525
rect 49145 3516 49157 3519
rect 49108 3488 49157 3516
rect 49108 3476 49114 3488
rect 49145 3485 49157 3488
rect 49191 3485 49203 3519
rect 49145 3479 49203 3485
rect 50525 3519 50583 3525
rect 50525 3485 50537 3519
rect 50571 3516 50583 3519
rect 50614 3516 50620 3528
rect 50571 3488 50620 3516
rect 50571 3485 50583 3488
rect 50525 3479 50583 3485
rect 50614 3476 50620 3488
rect 50672 3476 50678 3528
rect 50982 3476 50988 3528
rect 51040 3516 51046 3528
rect 51169 3519 51227 3525
rect 51169 3516 51181 3519
rect 51040 3488 51181 3516
rect 51040 3476 51046 3488
rect 51169 3485 51181 3488
rect 51215 3485 51227 3519
rect 51169 3479 51227 3485
rect 51534 3476 51540 3528
rect 51592 3516 51598 3528
rect 51813 3519 51871 3525
rect 51813 3516 51825 3519
rect 51592 3488 51825 3516
rect 51592 3476 51598 3488
rect 51813 3485 51825 3488
rect 51859 3485 51871 3519
rect 51813 3479 51871 3485
rect 46348 3420 47164 3448
rect 46348 3408 46354 3420
rect 23983 3352 26234 3380
rect 23983 3349 23995 3352
rect 23937 3343 23995 3349
rect 36354 3340 36360 3392
rect 36412 3380 36418 3392
rect 40034 3380 40040 3392
rect 36412 3352 40040 3380
rect 36412 3340 36418 3352
rect 40034 3340 40040 3352
rect 40092 3340 40098 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 24026 3176 24032 3188
rect 21468 3148 24032 3176
rect 21468 3049 21496 3148
rect 24026 3136 24032 3148
rect 24084 3136 24090 3188
rect 25774 3176 25780 3188
rect 24136 3148 25780 3176
rect 23934 3108 23940 3120
rect 22388 3080 23940 3108
rect 22388 3049 22416 3080
rect 23934 3068 23940 3080
rect 23992 3068 23998 3120
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21453 3043 21511 3049
rect 20855 3012 21404 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2972 13783 2975
rect 14366 2972 14372 2984
rect 13771 2944 14372 2972
rect 13771 2941 13783 2944
rect 13725 2935 13783 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 15657 2975 15715 2981
rect 15657 2941 15669 2975
rect 15703 2972 15715 2975
rect 16298 2972 16304 2984
rect 15703 2944 16304 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 19521 2975 19579 2981
rect 19521 2941 19533 2975
rect 19567 2972 19579 2975
rect 20898 2972 20904 2984
rect 19567 2944 20904 2972
rect 19567 2941 19579 2944
rect 19521 2935 19579 2941
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 21376 2972 21404 3012
rect 21453 3009 21465 3043
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 22373 3043 22431 3049
rect 22373 3009 22385 3043
rect 22419 3009 22431 3043
rect 22373 3003 22431 3009
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3040 22891 3043
rect 23290 3040 23296 3052
rect 22879 3012 23296 3040
rect 22879 3009 22891 3012
rect 22833 3003 22891 3009
rect 23290 3000 23296 3012
rect 23348 3000 23354 3052
rect 23750 3040 23756 3052
rect 23400 3012 23756 3040
rect 23400 2972 23428 3012
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 24026 3000 24032 3052
rect 24084 3040 24090 3052
rect 24136 3049 24164 3148
rect 25774 3136 25780 3148
rect 25832 3136 25838 3188
rect 36906 3136 36912 3188
rect 36964 3176 36970 3188
rect 36964 3148 39436 3176
rect 36964 3136 36970 3148
rect 24213 3111 24271 3117
rect 24213 3077 24225 3111
rect 24259 3108 24271 3111
rect 28994 3108 29000 3120
rect 24259 3080 29000 3108
rect 24259 3077 24271 3080
rect 24213 3071 24271 3077
rect 28994 3068 29000 3080
rect 29052 3068 29058 3120
rect 33965 3111 34023 3117
rect 33965 3077 33977 3111
rect 34011 3108 34023 3111
rect 34790 3108 34796 3120
rect 34011 3080 34796 3108
rect 34011 3077 34023 3080
rect 33965 3071 34023 3077
rect 34790 3068 34796 3080
rect 34848 3068 34854 3120
rect 36265 3111 36323 3117
rect 36265 3077 36277 3111
rect 36311 3108 36323 3111
rect 38197 3111 38255 3117
rect 38197 3108 38209 3111
rect 36311 3080 38209 3108
rect 36311 3077 36323 3080
rect 36265 3071 36323 3077
rect 38197 3077 38209 3080
rect 38243 3077 38255 3111
rect 38197 3071 38255 3077
rect 24121 3043 24179 3049
rect 24121 3040 24133 3043
rect 24084 3012 24133 3040
rect 24084 3000 24090 3012
rect 24121 3009 24133 3012
rect 24167 3009 24179 3043
rect 24121 3003 24179 3009
rect 24302 3000 24308 3052
rect 24360 3040 24366 3052
rect 24578 3040 24584 3052
rect 24360 3012 24584 3040
rect 24360 3000 24366 3012
rect 24578 3000 24584 3012
rect 24636 3000 24642 3052
rect 24762 3040 24768 3052
rect 24723 3012 24768 3040
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 34149 3043 34207 3049
rect 34149 3009 34161 3043
rect 34195 3040 34207 3043
rect 34698 3040 34704 3052
rect 34195 3012 34704 3040
rect 34195 3009 34207 3012
rect 34149 3003 34207 3009
rect 34698 3000 34704 3012
rect 34756 3000 34762 3052
rect 37366 3000 37372 3052
rect 37424 3040 37430 3052
rect 39408 3049 39436 3148
rect 37645 3043 37703 3049
rect 37645 3040 37657 3043
rect 37424 3012 37657 3040
rect 37424 3000 37430 3012
rect 37645 3009 37657 3012
rect 37691 3040 37703 3043
rect 38105 3043 38163 3049
rect 38105 3040 38117 3043
rect 37691 3012 38117 3040
rect 37691 3009 37703 3012
rect 37645 3003 37703 3009
rect 38105 3009 38117 3012
rect 38151 3009 38163 3043
rect 38105 3003 38163 3009
rect 39393 3043 39451 3049
rect 39393 3009 39405 3043
rect 39439 3009 39451 3043
rect 39393 3003 39451 3009
rect 42702 3000 42708 3052
rect 42760 3040 42766 3052
rect 43901 3043 43959 3049
rect 43901 3040 43913 3043
rect 42760 3012 43913 3040
rect 42760 3000 42766 3012
rect 43901 3009 43913 3012
rect 43947 3009 43959 3043
rect 43901 3003 43959 3009
rect 21376 2944 23428 2972
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 24949 2975 25007 2981
rect 24949 2972 24961 2975
rect 23532 2944 24961 2972
rect 23532 2932 23538 2944
rect 24949 2941 24961 2944
rect 24995 2941 25007 2975
rect 24949 2935 25007 2941
rect 26605 2975 26663 2981
rect 26605 2941 26617 2975
rect 26651 2972 26663 2975
rect 26970 2972 26976 2984
rect 26651 2944 26976 2972
rect 26651 2941 26663 2944
rect 26605 2935 26663 2941
rect 26970 2932 26976 2944
rect 27028 2932 27034 2984
rect 27617 2975 27675 2981
rect 27617 2941 27629 2975
rect 27663 2941 27675 2975
rect 27617 2935 27675 2941
rect 27801 2975 27859 2981
rect 27801 2941 27813 2975
rect 27847 2941 27859 2975
rect 29178 2972 29184 2984
rect 29139 2944 29184 2972
rect 27801 2935 27859 2941
rect 18877 2907 18935 2913
rect 18877 2873 18889 2907
rect 18923 2904 18935 2907
rect 20070 2904 20076 2916
rect 18923 2876 20076 2904
rect 18923 2873 18935 2876
rect 18877 2867 18935 2873
rect 20070 2864 20076 2876
rect 20128 2864 20134 2916
rect 20165 2907 20223 2913
rect 20165 2873 20177 2907
rect 20211 2904 20223 2907
rect 22554 2904 22560 2916
rect 20211 2876 22560 2904
rect 20211 2873 20223 2876
rect 20165 2867 20223 2873
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 23661 2907 23719 2913
rect 23661 2873 23673 2907
rect 23707 2904 23719 2907
rect 27632 2904 27660 2935
rect 23707 2876 27660 2904
rect 23707 2873 23719 2876
rect 23661 2867 23719 2873
rect 8202 2796 8208 2848
rect 8260 2836 8266 2848
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 8260 2808 8309 2836
rect 8260 2796 8266 2808
rect 8297 2805 8309 2808
rect 8343 2805 8355 2839
rect 8297 2799 8355 2805
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9674 2836 9680 2848
rect 9263 2808 9680 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9861 2839 9919 2845
rect 9861 2805 9873 2839
rect 9907 2836 9919 2839
rect 10226 2836 10232 2848
rect 9907 2808 10232 2836
rect 9907 2805 9919 2808
rect 9861 2799 9919 2805
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 10505 2839 10563 2845
rect 10505 2805 10517 2839
rect 10551 2836 10563 2839
rect 11054 2836 11060 2848
rect 10551 2808 11060 2836
rect 10551 2805 10563 2808
rect 10505 2799 10563 2805
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 11330 2836 11336 2848
rect 11195 2808 11336 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2836 12495 2839
rect 12710 2836 12716 2848
rect 12483 2808 12716 2836
rect 12483 2805 12495 2808
rect 12437 2799 12495 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13538 2836 13544 2848
rect 13127 2808 13544 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 14642 2836 14648 2848
rect 14415 2808 14648 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 15013 2839 15071 2845
rect 15013 2805 15025 2839
rect 15059 2836 15071 2839
rect 15470 2836 15476 2848
rect 15059 2808 15476 2836
rect 15059 2805 15071 2808
rect 15013 2799 15071 2805
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 16850 2836 16856 2848
rect 16347 2808 16856 2836
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 17589 2839 17647 2845
rect 17589 2805 17601 2839
rect 17635 2836 17647 2839
rect 18138 2836 18144 2848
rect 17635 2808 18144 2836
rect 17635 2805 17647 2808
rect 17589 2799 17647 2805
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 18233 2839 18291 2845
rect 18233 2805 18245 2839
rect 18279 2836 18291 2839
rect 18690 2836 18696 2848
rect 18279 2808 18696 2836
rect 18279 2805 18291 2808
rect 18233 2799 18291 2805
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 22925 2839 22983 2845
rect 22925 2805 22937 2839
rect 22971 2836 22983 2839
rect 24578 2836 24584 2848
rect 22971 2808 24584 2836
rect 22971 2805 22983 2808
rect 22925 2799 22983 2805
rect 24578 2796 24584 2808
rect 24636 2796 24642 2848
rect 24854 2796 24860 2848
rect 24912 2836 24918 2848
rect 27816 2836 27844 2935
rect 29178 2932 29184 2944
rect 29236 2932 29242 2984
rect 29917 2975 29975 2981
rect 29917 2941 29929 2975
rect 29963 2941 29975 2975
rect 30098 2972 30104 2984
rect 30059 2944 30104 2972
rect 29917 2935 29975 2941
rect 27890 2864 27896 2916
rect 27948 2904 27954 2916
rect 29932 2904 29960 2935
rect 30098 2932 30104 2944
rect 30156 2932 30162 2984
rect 31110 2972 31116 2984
rect 31071 2944 31116 2972
rect 31110 2932 31116 2944
rect 31168 2932 31174 2984
rect 31938 2932 31944 2984
rect 31996 2972 32002 2984
rect 32309 2975 32367 2981
rect 32309 2972 32321 2975
rect 31996 2944 32321 2972
rect 31996 2932 32002 2944
rect 32309 2941 32321 2944
rect 32355 2941 32367 2975
rect 32309 2935 32367 2941
rect 34422 2932 34428 2984
rect 34480 2972 34486 2984
rect 34609 2975 34667 2981
rect 34609 2972 34621 2975
rect 34480 2944 34621 2972
rect 34480 2932 34486 2944
rect 34609 2941 34621 2944
rect 34655 2941 34667 2975
rect 34609 2935 34667 2941
rect 36449 2975 36507 2981
rect 36449 2941 36461 2975
rect 36495 2972 36507 2975
rect 37458 2972 37464 2984
rect 36495 2944 37464 2972
rect 36495 2941 36507 2944
rect 36449 2935 36507 2941
rect 37458 2932 37464 2944
rect 37516 2932 37522 2984
rect 38749 2975 38807 2981
rect 38749 2972 38761 2975
rect 37568 2944 38761 2972
rect 27948 2876 29960 2904
rect 27948 2864 27954 2876
rect 36078 2864 36084 2916
rect 36136 2904 36142 2916
rect 37568 2904 37596 2944
rect 38749 2941 38761 2944
rect 38795 2941 38807 2975
rect 38749 2935 38807 2941
rect 38838 2932 38844 2984
rect 38896 2972 38902 2984
rect 40681 2975 40739 2981
rect 40681 2972 40693 2975
rect 38896 2944 40693 2972
rect 38896 2932 38902 2944
rect 40681 2941 40693 2944
rect 40727 2941 40739 2975
rect 40681 2935 40739 2941
rect 40770 2932 40776 2984
rect 40828 2972 40834 2984
rect 42613 2975 42671 2981
rect 42613 2972 42625 2975
rect 40828 2944 42625 2972
rect 40828 2932 40834 2944
rect 42613 2941 42625 2944
rect 42659 2941 42671 2975
rect 42613 2935 42671 2941
rect 43254 2932 43260 2984
rect 43312 2972 43318 2984
rect 44545 2975 44603 2981
rect 44545 2972 44557 2975
rect 43312 2944 44557 2972
rect 43312 2932 43318 2944
rect 44545 2941 44557 2944
rect 44591 2941 44603 2975
rect 45833 2975 45891 2981
rect 45833 2972 45845 2975
rect 44545 2935 44603 2941
rect 45526 2944 45845 2972
rect 36136 2876 37596 2904
rect 36136 2864 36142 2876
rect 37734 2864 37740 2916
rect 37792 2904 37798 2916
rect 37792 2876 39528 2904
rect 37792 2864 37798 2876
rect 24912 2808 27844 2836
rect 24912 2796 24918 2808
rect 29454 2796 29460 2848
rect 29512 2836 29518 2848
rect 30190 2836 30196 2848
rect 29512 2808 30196 2836
rect 29512 2796 29518 2808
rect 30190 2796 30196 2808
rect 30248 2796 30254 2848
rect 37550 2836 37556 2848
rect 37511 2808 37556 2836
rect 37550 2796 37556 2808
rect 37608 2796 37614 2848
rect 39500 2836 39528 2876
rect 39666 2864 39672 2916
rect 39724 2904 39730 2916
rect 41325 2907 41383 2913
rect 41325 2904 41337 2907
rect 39724 2876 41337 2904
rect 39724 2864 39730 2876
rect 41325 2873 41337 2876
rect 41371 2873 41383 2907
rect 41325 2867 41383 2873
rect 41598 2864 41604 2916
rect 41656 2904 41662 2916
rect 41656 2876 42748 2904
rect 41656 2864 41662 2876
rect 40037 2839 40095 2845
rect 40037 2836 40049 2839
rect 39500 2808 40049 2836
rect 40037 2805 40049 2808
rect 40083 2805 40095 2839
rect 42720 2836 42748 2876
rect 44910 2864 44916 2916
rect 44968 2904 44974 2916
rect 45526 2904 45554 2944
rect 45833 2941 45845 2944
rect 45879 2941 45891 2975
rect 45833 2935 45891 2941
rect 48774 2932 48780 2984
rect 48832 2972 48838 2984
rect 49697 2975 49755 2981
rect 49697 2972 49709 2975
rect 48832 2944 49709 2972
rect 48832 2932 48838 2944
rect 49697 2941 49709 2944
rect 49743 2941 49755 2975
rect 49697 2935 49755 2941
rect 46477 2907 46535 2913
rect 46477 2904 46489 2907
rect 44968 2876 45554 2904
rect 45756 2876 46489 2904
rect 44968 2864 44974 2876
rect 43257 2839 43315 2845
rect 43257 2836 43269 2839
rect 42720 2808 43269 2836
rect 40037 2799 40095 2805
rect 43257 2805 43269 2808
rect 43303 2805 43315 2839
rect 43257 2799 43315 2805
rect 43806 2796 43812 2848
rect 43864 2836 43870 2848
rect 45189 2839 45247 2845
rect 45189 2836 45201 2839
rect 43864 2808 45201 2836
rect 43864 2796 43870 2808
rect 45189 2805 45201 2808
rect 45235 2805 45247 2839
rect 45189 2799 45247 2805
rect 45462 2796 45468 2848
rect 45520 2836 45526 2848
rect 45756 2836 45784 2876
rect 46477 2873 46489 2876
rect 46523 2873 46535 2907
rect 46477 2867 46535 2873
rect 47670 2864 47676 2916
rect 47728 2904 47734 2916
rect 48409 2907 48467 2913
rect 48409 2904 48421 2907
rect 47728 2876 48421 2904
rect 47728 2864 47734 2876
rect 48409 2873 48421 2876
rect 48455 2873 48467 2907
rect 48409 2867 48467 2873
rect 49602 2864 49608 2916
rect 49660 2904 49666 2916
rect 50341 2907 50399 2913
rect 50341 2904 50353 2907
rect 49660 2876 50353 2904
rect 49660 2864 49666 2876
rect 50341 2873 50353 2876
rect 50387 2873 50399 2907
rect 50341 2867 50399 2873
rect 50706 2864 50712 2916
rect 50764 2904 50770 2916
rect 51629 2907 51687 2913
rect 51629 2904 51641 2907
rect 50764 2876 51641 2904
rect 50764 2864 50770 2876
rect 51629 2873 51641 2876
rect 51675 2873 51687 2907
rect 51629 2867 51687 2873
rect 45520 2808 45784 2836
rect 45520 2796 45526 2808
rect 46842 2796 46848 2848
rect 46900 2836 46906 2848
rect 47765 2839 47823 2845
rect 47765 2836 47777 2839
rect 46900 2808 47777 2836
rect 46900 2796 46906 2808
rect 47765 2805 47777 2808
rect 47811 2805 47823 2839
rect 47765 2799 47823 2805
rect 48222 2796 48228 2848
rect 48280 2836 48286 2848
rect 49053 2839 49111 2845
rect 49053 2836 49065 2839
rect 48280 2808 49065 2836
rect 48280 2796 48286 2808
rect 49053 2805 49065 2808
rect 49099 2805 49111 2839
rect 49053 2799 49111 2805
rect 50154 2796 50160 2848
rect 50212 2836 50218 2848
rect 50985 2839 51043 2845
rect 50985 2836 50997 2839
rect 50212 2808 50997 2836
rect 50212 2796 50218 2808
rect 50985 2805 50997 2808
rect 51031 2805 51043 2839
rect 50985 2799 51043 2805
rect 52086 2796 52092 2848
rect 52144 2836 52150 2848
rect 52917 2839 52975 2845
rect 52917 2836 52929 2839
rect 52144 2808 52929 2836
rect 52144 2796 52150 2808
rect 52917 2805 52929 2808
rect 52963 2805 52975 2839
rect 52917 2799 52975 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 23293 2635 23351 2641
rect 23293 2601 23305 2635
rect 23339 2632 23351 2635
rect 23474 2632 23480 2644
rect 23339 2604 23480 2632
rect 23339 2601 23351 2604
rect 23293 2595 23351 2601
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 23937 2635 23995 2641
rect 23937 2601 23949 2635
rect 23983 2632 23995 2635
rect 24854 2632 24860 2644
rect 23983 2604 24860 2632
rect 23983 2601 23995 2604
rect 23937 2595 23995 2601
rect 24854 2592 24860 2604
rect 24912 2592 24918 2644
rect 26206 2604 29776 2632
rect 7929 2567 7987 2573
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 8570 2564 8576 2576
rect 7975 2536 8576 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 8570 2524 8576 2536
rect 8628 2524 8634 2576
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 10502 2564 10508 2576
rect 9907 2536 10508 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 13725 2567 13783 2573
rect 13725 2533 13737 2567
rect 13771 2564 13783 2567
rect 15194 2564 15200 2576
rect 13771 2536 15200 2564
rect 13771 2533 13783 2536
rect 13725 2527 13783 2533
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 15657 2567 15715 2573
rect 15657 2533 15669 2567
rect 15703 2564 15715 2567
rect 17126 2564 17132 2576
rect 15703 2536 17132 2564
rect 15703 2533 15715 2536
rect 15657 2527 15715 2533
rect 17126 2524 17132 2536
rect 17184 2524 17190 2576
rect 17589 2567 17647 2573
rect 17589 2533 17601 2567
rect 17635 2564 17647 2567
rect 18966 2564 18972 2576
rect 17635 2536 18972 2564
rect 17635 2533 17647 2536
rect 17589 2527 17647 2533
rect 18966 2524 18972 2536
rect 19024 2524 19030 2576
rect 22649 2567 22707 2573
rect 22649 2533 22661 2567
rect 22695 2564 22707 2567
rect 23566 2564 23572 2576
rect 22695 2536 23572 2564
rect 22695 2533 22707 2536
rect 22649 2527 22707 2533
rect 23566 2524 23572 2536
rect 23624 2524 23630 2576
rect 25317 2567 25375 2573
rect 25317 2533 25329 2567
rect 25363 2564 25375 2567
rect 26206 2564 26234 2604
rect 25363 2536 26234 2564
rect 26436 2536 27568 2564
rect 25363 2533 25375 2536
rect 25317 2527 25375 2533
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 13814 2496 13820 2508
rect 13127 2468 13820 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 13814 2456 13820 2468
rect 13872 2456 13878 2508
rect 16301 2499 16359 2505
rect 16301 2465 16313 2499
rect 16347 2496 16359 2499
rect 17862 2496 17868 2508
rect 16347 2468 17868 2496
rect 16347 2465 16359 2468
rect 16301 2459 16359 2465
rect 17862 2456 17868 2468
rect 17920 2456 17926 2508
rect 18233 2499 18291 2505
rect 18233 2465 18245 2499
rect 18279 2496 18291 2499
rect 19978 2496 19984 2508
rect 18279 2468 19984 2496
rect 18279 2465 18291 2468
rect 18233 2459 18291 2465
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 20165 2499 20223 2505
rect 20165 2465 20177 2499
rect 20211 2496 20223 2499
rect 23382 2496 23388 2508
rect 20211 2468 23388 2496
rect 20211 2465 20223 2468
rect 20165 2459 20223 2465
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 24578 2456 24584 2508
rect 24636 2496 24642 2508
rect 26436 2496 26464 2536
rect 27540 2505 27568 2536
rect 27341 2499 27399 2505
rect 27341 2496 27353 2499
rect 24636 2468 26464 2496
rect 26528 2468 27353 2496
rect 24636 2456 24642 2468
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7650 2428 7656 2440
rect 7331 2400 7656 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2428 8631 2431
rect 9306 2428 9312 2440
rect 8619 2400 9312 2428
rect 8619 2397 8631 2400
rect 8573 2391 8631 2397
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2428 11207 2431
rect 12158 2428 12164 2440
rect 11195 2400 12164 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 10520 2360 10548 2391
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12986 2428 12992 2440
rect 12483 2400 12992 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 16022 2428 16028 2440
rect 15059 2400 16028 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2428 20867 2431
rect 21453 2431 21511 2437
rect 20855 2400 21404 2428
rect 20855 2397 20867 2400
rect 20809 2391 20867 2397
rect 11882 2360 11888 2372
rect 10520 2332 11888 2360
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 18892 2360 18920 2391
rect 21174 2360 21180 2372
rect 18892 2332 21180 2360
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 21376 2292 21404 2400
rect 21453 2397 21465 2431
rect 21499 2397 21511 2431
rect 21453 2391 21511 2397
rect 22741 2431 22799 2437
rect 22741 2397 22753 2431
rect 22787 2428 22799 2431
rect 23201 2431 23259 2437
rect 23201 2428 23213 2431
rect 22787 2400 23213 2428
rect 22787 2397 22799 2400
rect 22741 2391 22799 2397
rect 23201 2397 23213 2400
rect 23247 2428 23259 2431
rect 23290 2428 23296 2440
rect 23247 2400 23296 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 21468 2360 21496 2391
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 24026 2428 24032 2440
rect 23987 2400 24032 2428
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 25774 2428 25780 2440
rect 25735 2400 25780 2428
rect 25774 2388 25780 2400
rect 25832 2388 25838 2440
rect 25866 2388 25872 2440
rect 25924 2428 25930 2440
rect 26528 2428 26556 2468
rect 27341 2465 27353 2468
rect 27387 2465 27399 2499
rect 27341 2459 27399 2465
rect 27525 2499 27583 2505
rect 27525 2465 27537 2499
rect 27571 2465 27583 2499
rect 28534 2496 28540 2508
rect 28495 2468 28540 2496
rect 27525 2459 27583 2465
rect 28534 2456 28540 2468
rect 28592 2456 28598 2508
rect 29748 2505 29776 2604
rect 34606 2592 34612 2644
rect 34664 2632 34670 2644
rect 34977 2635 35035 2641
rect 34977 2632 34989 2635
rect 34664 2604 34989 2632
rect 34664 2592 34670 2604
rect 34977 2601 34989 2604
rect 35023 2601 35035 2635
rect 37458 2632 37464 2644
rect 37419 2604 37464 2632
rect 34977 2595 35035 2601
rect 37458 2592 37464 2604
rect 37516 2592 37522 2644
rect 38746 2632 38752 2644
rect 38707 2604 38752 2632
rect 38746 2592 38752 2604
rect 38804 2592 38810 2644
rect 40034 2632 40040 2644
rect 39995 2604 40040 2632
rect 40034 2592 40040 2604
rect 40092 2592 40098 2644
rect 34698 2524 34704 2576
rect 34756 2564 34762 2576
rect 35529 2567 35587 2573
rect 35529 2564 35541 2567
rect 34756 2536 35541 2564
rect 34756 2524 34762 2536
rect 35529 2533 35541 2536
rect 35575 2533 35587 2567
rect 35529 2527 35587 2533
rect 42150 2524 42156 2576
rect 42208 2564 42214 2576
rect 43901 2567 43959 2573
rect 43901 2564 43913 2567
rect 42208 2536 43913 2564
rect 42208 2524 42214 2536
rect 43901 2533 43913 2536
rect 43947 2533 43959 2567
rect 43901 2527 43959 2533
rect 44634 2524 44640 2576
rect 44692 2564 44698 2576
rect 46477 2567 46535 2573
rect 46477 2564 46489 2567
rect 44692 2536 46489 2564
rect 44692 2524 44698 2536
rect 46477 2533 46489 2536
rect 46523 2533 46535 2567
rect 46477 2527 46535 2533
rect 48498 2524 48504 2576
rect 48556 2564 48562 2576
rect 50341 2567 50399 2573
rect 50341 2564 50353 2567
rect 48556 2536 50353 2564
rect 48556 2524 48562 2536
rect 50341 2533 50353 2536
rect 50387 2533 50399 2567
rect 50341 2527 50399 2533
rect 51810 2524 51816 2576
rect 51868 2564 51874 2576
rect 53561 2567 53619 2573
rect 53561 2564 53573 2567
rect 51868 2536 53573 2564
rect 51868 2524 51874 2536
rect 53561 2533 53573 2536
rect 53607 2533 53619 2567
rect 53561 2527 53619 2533
rect 29733 2499 29791 2505
rect 29733 2465 29745 2499
rect 29779 2465 29791 2499
rect 30190 2496 30196 2508
rect 30151 2468 30196 2496
rect 29733 2459 29791 2465
rect 30190 2456 30196 2468
rect 30248 2456 30254 2508
rect 33318 2496 33324 2508
rect 33279 2468 33324 2496
rect 33318 2456 33324 2468
rect 33376 2456 33382 2508
rect 34333 2499 34391 2505
rect 34333 2465 34345 2499
rect 34379 2496 34391 2499
rect 35434 2496 35440 2508
rect 34379 2468 35440 2496
rect 34379 2465 34391 2468
rect 34333 2459 34391 2465
rect 35434 2456 35440 2468
rect 35492 2456 35498 2508
rect 38010 2456 38016 2508
rect 38068 2496 38074 2508
rect 40681 2499 40739 2505
rect 40681 2496 40693 2499
rect 38068 2468 40693 2496
rect 38068 2456 38074 2468
rect 40681 2465 40693 2468
rect 40727 2465 40739 2499
rect 40681 2459 40739 2465
rect 41414 2456 41420 2508
rect 41472 2496 41478 2508
rect 43257 2499 43315 2505
rect 43257 2496 43269 2499
rect 41472 2468 43269 2496
rect 41472 2456 41478 2468
rect 43257 2465 43269 2468
rect 43303 2465 43315 2499
rect 43257 2459 43315 2465
rect 43530 2456 43536 2508
rect 43588 2496 43594 2508
rect 45189 2499 45247 2505
rect 45189 2496 45201 2499
rect 43588 2468 45201 2496
rect 43588 2456 43594 2468
rect 45189 2465 45201 2468
rect 45235 2465 45247 2499
rect 45189 2459 45247 2465
rect 46566 2456 46572 2508
rect 46624 2496 46630 2508
rect 48409 2499 48467 2505
rect 48409 2496 48421 2499
rect 46624 2468 48421 2496
rect 46624 2456 46630 2468
rect 48409 2465 48421 2468
rect 48455 2465 48467 2499
rect 48409 2459 48467 2465
rect 49326 2456 49332 2508
rect 49384 2496 49390 2508
rect 50985 2499 51043 2505
rect 50985 2496 50997 2499
rect 49384 2468 50997 2496
rect 49384 2456 49390 2468
rect 50985 2465 50997 2468
rect 51031 2465 51043 2499
rect 50985 2459 51043 2465
rect 52362 2456 52368 2508
rect 52420 2496 52426 2508
rect 54205 2499 54263 2505
rect 54205 2496 54217 2499
rect 52420 2468 54217 2496
rect 52420 2456 52426 2468
rect 54205 2465 54217 2468
rect 54251 2465 54263 2499
rect 54205 2459 54263 2465
rect 25924 2400 26556 2428
rect 26605 2431 26663 2437
rect 25924 2388 25930 2400
rect 26605 2397 26617 2431
rect 26651 2397 26663 2431
rect 26605 2391 26663 2397
rect 35069 2431 35127 2437
rect 35069 2397 35081 2431
rect 35115 2428 35127 2431
rect 35618 2428 35624 2440
rect 35115 2400 35624 2428
rect 35115 2397 35127 2400
rect 35069 2391 35127 2397
rect 25590 2360 25596 2372
rect 21468 2332 25596 2360
rect 25590 2320 25596 2332
rect 25648 2320 25654 2372
rect 26620 2360 26648 2391
rect 35618 2388 35624 2400
rect 35676 2428 35682 2440
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 35676 2400 36369 2428
rect 35676 2388 35682 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 38105 2431 38163 2437
rect 38105 2397 38117 2431
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 27890 2360 27896 2372
rect 26620 2332 27896 2360
rect 27890 2320 27896 2332
rect 27948 2320 27954 2372
rect 28994 2320 29000 2372
rect 29052 2360 29058 2372
rect 29917 2363 29975 2369
rect 29917 2360 29929 2363
rect 29052 2332 29929 2360
rect 29052 2320 29058 2332
rect 29917 2329 29929 2332
rect 29963 2329 29975 2363
rect 29917 2323 29975 2329
rect 34149 2363 34207 2369
rect 34149 2329 34161 2363
rect 34195 2360 34207 2363
rect 34698 2360 34704 2372
rect 34195 2332 34704 2360
rect 34195 2329 34207 2332
rect 34149 2323 34207 2329
rect 34698 2320 34704 2332
rect 34756 2320 34762 2372
rect 34790 2320 34796 2372
rect 34848 2360 34854 2372
rect 36265 2363 36323 2369
rect 36265 2360 36277 2363
rect 34848 2332 36277 2360
rect 34848 2320 34854 2332
rect 36265 2329 36277 2332
rect 36311 2329 36323 2363
rect 36265 2323 36323 2329
rect 25038 2292 25044 2304
rect 21376 2264 25044 2292
rect 25038 2252 25044 2264
rect 25096 2252 25102 2304
rect 25869 2295 25927 2301
rect 25869 2261 25881 2295
rect 25915 2292 25927 2295
rect 30098 2292 30104 2304
rect 25915 2264 30104 2292
rect 25915 2261 25927 2264
rect 25869 2255 25927 2261
rect 30098 2252 30104 2264
rect 30156 2252 30162 2304
rect 34974 2252 34980 2304
rect 35032 2292 35038 2304
rect 38120 2292 38148 2391
rect 38562 2388 38568 2440
rect 38620 2428 38626 2440
rect 41325 2431 41383 2437
rect 41325 2428 41337 2431
rect 38620 2400 41337 2428
rect 38620 2388 38626 2400
rect 41325 2397 41337 2400
rect 41371 2397 41383 2431
rect 41325 2391 41383 2397
rect 42613 2431 42671 2437
rect 42613 2397 42625 2431
rect 42659 2397 42671 2431
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 42613 2391 42671 2397
rect 45526 2400 45845 2428
rect 40218 2320 40224 2372
rect 40276 2360 40282 2372
rect 42628 2360 42656 2391
rect 40276 2332 42656 2360
rect 40276 2320 40282 2332
rect 44082 2320 44088 2372
rect 44140 2360 44146 2372
rect 45526 2360 45554 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 45833 2391 45891 2397
rect 46014 2388 46020 2440
rect 46072 2428 46078 2440
rect 47765 2431 47823 2437
rect 47765 2428 47777 2431
rect 46072 2400 47777 2428
rect 46072 2388 46078 2400
rect 47765 2397 47777 2400
rect 47811 2397 47823 2431
rect 47765 2391 47823 2397
rect 49053 2431 49111 2437
rect 49053 2397 49065 2431
rect 49099 2397 49111 2431
rect 49053 2391 49111 2397
rect 44140 2332 45554 2360
rect 44140 2320 44146 2332
rect 47394 2320 47400 2372
rect 47452 2360 47458 2372
rect 49068 2360 49096 2391
rect 49878 2388 49884 2440
rect 49936 2428 49942 2440
rect 51629 2431 51687 2437
rect 51629 2428 51641 2431
rect 49936 2400 51641 2428
rect 49936 2388 49942 2400
rect 51629 2397 51641 2400
rect 51675 2397 51687 2431
rect 51629 2391 51687 2397
rect 52917 2431 52975 2437
rect 52917 2397 52929 2431
rect 52963 2397 52975 2431
rect 52917 2391 52975 2397
rect 47452 2332 49096 2360
rect 47452 2320 47458 2332
rect 51258 2320 51264 2372
rect 51316 2360 51322 2372
rect 52932 2360 52960 2391
rect 51316 2332 52960 2360
rect 51316 2320 51322 2332
rect 35032 2264 38148 2292
rect 35032 2252 35038 2264
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 34698 2048 34704 2100
rect 34756 2088 34762 2100
rect 37550 2088 37556 2100
rect 34756 2060 37556 2088
rect 34756 2048 34762 2060
rect 37550 2048 37556 2060
rect 37608 2048 37614 2100
rect 23750 1436 23756 1488
rect 23808 1476 23814 1488
rect 24210 1476 24216 1488
rect 23808 1448 24216 1476
rect 23808 1436 23814 1448
rect 24210 1436 24216 1448
rect 24268 1436 24274 1488
rect 34698 1368 34704 1420
rect 34756 1408 34762 1420
rect 35710 1408 35716 1420
rect 34756 1380 35716 1408
rect 34756 1368 34762 1380
rect 35710 1368 35716 1380
rect 35768 1368 35774 1420
<< via1 >>
rect 21364 57876 21416 57928
rect 27436 57876 27488 57928
rect 33416 57876 33468 57928
rect 17868 57808 17920 57860
rect 28448 57808 28500 57860
rect 22836 57740 22888 57792
rect 23940 57740 23992 57792
rect 24768 57740 24820 57792
rect 30564 57808 30616 57860
rect 41420 57808 41472 57860
rect 45928 57808 45980 57860
rect 29184 57740 29236 57792
rect 33968 57740 34020 57792
rect 42892 57740 42944 57792
rect 46848 57740 46900 57792
rect 54116 57740 54168 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 3700 57536 3752 57588
rect 5080 57536 5132 57588
rect 10600 57536 10652 57588
rect 11980 57536 12032 57588
rect 13360 57536 13412 57588
rect 14740 57536 14792 57588
rect 16120 57536 16172 57588
rect 17500 57536 17552 57588
rect 19340 57536 19392 57588
rect 20260 57536 20312 57588
rect 22192 57536 22244 57588
rect 23020 57536 23072 57588
rect 25044 57536 25096 57588
rect 25780 57536 25832 57588
rect 27160 57536 27212 57588
rect 28540 57536 28592 57588
rect 7380 57400 7432 57452
rect 7840 57400 7892 57452
rect 8760 57400 8812 57452
rect 9220 57400 9272 57452
rect 10140 57400 10192 57452
rect 10968 57443 11020 57452
rect 10968 57409 10977 57443
rect 10977 57409 11011 57443
rect 11011 57409 11020 57443
rect 10968 57400 11020 57409
rect 12348 57443 12400 57452
rect 12348 57409 12357 57443
rect 12357 57409 12391 57443
rect 12391 57409 12400 57443
rect 12348 57400 12400 57409
rect 12900 57400 12952 57452
rect 6092 57332 6144 57384
rect 5448 57264 5500 57316
rect 15660 57400 15712 57452
rect 17132 57443 17184 57452
rect 17132 57409 17141 57443
rect 17141 57409 17175 57443
rect 17175 57409 17184 57443
rect 17132 57400 17184 57409
rect 17868 57443 17920 57452
rect 17868 57409 17877 57443
rect 17877 57409 17911 57443
rect 17911 57409 17920 57443
rect 17868 57400 17920 57409
rect 18420 57400 18472 57452
rect 23480 57468 23532 57520
rect 24400 57468 24452 57520
rect 23204 57443 23256 57452
rect 22744 57332 22796 57384
rect 23204 57409 23213 57443
rect 23213 57409 23247 57443
rect 23247 57409 23256 57443
rect 23204 57400 23256 57409
rect 23664 57443 23716 57452
rect 23664 57409 23673 57443
rect 23673 57409 23707 57443
rect 23707 57409 23716 57443
rect 23664 57400 23716 57409
rect 23756 57400 23808 57452
rect 24768 57443 24820 57452
rect 24768 57409 24777 57443
rect 24777 57409 24811 57443
rect 24811 57409 24820 57443
rect 24768 57400 24820 57409
rect 29184 57468 29236 57520
rect 25136 57400 25188 57452
rect 27252 57443 27304 57452
rect 27252 57409 27261 57443
rect 27261 57409 27295 57443
rect 27295 57409 27304 57443
rect 27252 57400 27304 57409
rect 25228 57332 25280 57384
rect 22836 57196 22888 57248
rect 23480 57264 23532 57316
rect 23572 57264 23624 57316
rect 29276 57400 29328 57452
rect 31576 57468 31628 57520
rect 34520 57536 34572 57588
rect 45744 57536 45796 57588
rect 54116 57536 54168 57588
rect 34244 57468 34296 57520
rect 30472 57400 30524 57452
rect 30840 57443 30892 57452
rect 30840 57409 30849 57443
rect 30849 57409 30883 57443
rect 30883 57409 30892 57443
rect 30840 57400 30892 57409
rect 30012 57332 30064 57384
rect 30288 57264 30340 57316
rect 31852 57332 31904 57384
rect 32036 57332 32088 57384
rect 32588 57375 32640 57384
rect 32588 57341 32597 57375
rect 32597 57341 32631 57375
rect 32631 57341 32640 57375
rect 32588 57332 32640 57341
rect 33508 57400 33560 57452
rect 34152 57400 34204 57452
rect 35532 57443 35584 57452
rect 34336 57332 34388 57384
rect 35532 57409 35541 57443
rect 35541 57409 35575 57443
rect 35575 57409 35584 57443
rect 35532 57400 35584 57409
rect 35900 57400 35952 57452
rect 37280 57400 37332 57452
rect 38660 57400 38712 57452
rect 39856 57400 39908 57452
rect 45560 57468 45612 57520
rect 41052 57400 41104 57452
rect 42800 57400 42852 57452
rect 44088 57400 44140 57452
rect 44272 57400 44324 57452
rect 44456 57400 44508 57452
rect 44916 57400 44968 57452
rect 47400 57400 47452 57452
rect 49700 57400 49752 57452
rect 52460 57468 52512 57520
rect 53012 57511 53064 57520
rect 53012 57477 53021 57511
rect 53021 57477 53055 57511
rect 53055 57477 53064 57511
rect 53012 57468 53064 57477
rect 51080 57400 51132 57452
rect 51448 57400 51500 57452
rect 53840 57400 53892 57452
rect 54300 57400 54352 57452
rect 55220 57400 55272 57452
rect 55772 57443 55824 57452
rect 55772 57409 55781 57443
rect 55781 57409 55815 57443
rect 55815 57409 55824 57443
rect 55772 57400 55824 57409
rect 56140 57400 56192 57452
rect 35716 57332 35768 57384
rect 36268 57375 36320 57384
rect 36268 57341 36277 57375
rect 36277 57341 36311 57375
rect 36311 57341 36320 57375
rect 36268 57332 36320 57341
rect 36636 57332 36688 57384
rect 41788 57375 41840 57384
rect 41788 57341 41797 57375
rect 41797 57341 41831 57375
rect 41831 57341 41840 57375
rect 41788 57332 41840 57341
rect 42984 57332 43036 57384
rect 43628 57332 43680 57384
rect 43996 57332 44048 57384
rect 45744 57332 45796 57384
rect 46940 57332 46992 57384
rect 23848 57196 23900 57248
rect 24032 57239 24084 57248
rect 24032 57205 24041 57239
rect 24041 57205 24075 57239
rect 24075 57205 24084 57239
rect 24032 57196 24084 57205
rect 24124 57196 24176 57248
rect 25320 57196 25372 57248
rect 28816 57196 28868 57248
rect 28908 57196 28960 57248
rect 36728 57264 36780 57316
rect 38936 57264 38988 57316
rect 40684 57264 40736 57316
rect 41236 57264 41288 57316
rect 45652 57264 45704 57316
rect 55680 57332 55732 57384
rect 31576 57196 31628 57248
rect 38752 57239 38804 57248
rect 38752 57205 38761 57239
rect 38761 57205 38795 57239
rect 38795 57205 38804 57239
rect 38752 57196 38804 57205
rect 40500 57196 40552 57248
rect 43352 57196 43404 57248
rect 45468 57196 45520 57248
rect 46388 57239 46440 57248
rect 46388 57205 46397 57239
rect 46397 57205 46431 57239
rect 46431 57205 46440 57239
rect 46388 57196 46440 57205
rect 47032 57239 47084 57248
rect 47032 57205 47041 57239
rect 47041 57205 47075 57239
rect 47075 57205 47084 57239
rect 47032 57196 47084 57205
rect 51816 57239 51868 57248
rect 51816 57205 51825 57239
rect 51825 57205 51859 57239
rect 51859 57205 51868 57239
rect 51816 57196 51868 57205
rect 53104 57239 53156 57248
rect 53104 57205 53113 57239
rect 53113 57205 53147 57239
rect 53147 57205 53156 57239
rect 53104 57196 53156 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 4620 56992 4672 57044
rect 6000 56992 6052 57044
rect 6460 56992 6512 57044
rect 11520 56992 11572 57044
rect 14280 56992 14332 57044
rect 17040 56992 17092 57044
rect 19984 56992 20036 57044
rect 21180 56992 21232 57044
rect 21640 56992 21692 57044
rect 23204 56992 23256 57044
rect 23848 56992 23900 57044
rect 27160 56992 27212 57044
rect 27436 56992 27488 57044
rect 27620 56992 27672 57044
rect 28908 56992 28960 57044
rect 31300 57035 31352 57044
rect 31300 57001 31309 57035
rect 31309 57001 31343 57035
rect 31343 57001 31352 57035
rect 31300 56992 31352 57001
rect 10968 56924 11020 56976
rect 21364 56924 21416 56976
rect 24124 56924 24176 56976
rect 22744 56856 22796 56908
rect 23756 56856 23808 56908
rect 25044 56899 25096 56908
rect 25044 56865 25053 56899
rect 25053 56865 25087 56899
rect 25087 56865 25096 56899
rect 25044 56856 25096 56865
rect 23480 56788 23532 56840
rect 24768 56788 24820 56840
rect 25136 56831 25188 56840
rect 25136 56797 25145 56831
rect 25145 56797 25179 56831
rect 25179 56797 25188 56831
rect 25136 56788 25188 56797
rect 25688 56788 25740 56840
rect 28356 56924 28408 56976
rect 28448 56924 28500 56976
rect 28816 56967 28868 56976
rect 28816 56933 28825 56967
rect 28825 56933 28859 56967
rect 28859 56933 28868 56967
rect 28816 56924 28868 56933
rect 36452 56992 36504 57044
rect 36544 56992 36596 57044
rect 41052 57035 41104 57044
rect 28264 56856 28316 56908
rect 27436 56831 27488 56840
rect 27436 56797 27445 56831
rect 27445 56797 27479 56831
rect 27479 56797 27488 56831
rect 27436 56788 27488 56797
rect 27528 56831 27580 56840
rect 27528 56797 27537 56831
rect 27537 56797 27571 56831
rect 27571 56797 27580 56831
rect 27804 56831 27856 56840
rect 27528 56788 27580 56797
rect 27804 56797 27813 56831
rect 27813 56797 27847 56831
rect 27847 56797 27856 56831
rect 27804 56788 27856 56797
rect 22192 56720 22244 56772
rect 23848 56695 23900 56704
rect 23848 56661 23857 56695
rect 23857 56661 23891 56695
rect 23891 56661 23900 56695
rect 23848 56652 23900 56661
rect 25596 56652 25648 56704
rect 27528 56652 27580 56704
rect 28724 56652 28776 56704
rect 29276 56856 29328 56908
rect 30012 56856 30064 56908
rect 31944 56924 31996 56976
rect 33968 56924 34020 56976
rect 29184 56831 29236 56840
rect 29184 56797 29193 56831
rect 29193 56797 29227 56831
rect 29227 56797 29236 56831
rect 29184 56788 29236 56797
rect 30288 56831 30340 56840
rect 30012 56720 30064 56772
rect 30288 56797 30297 56831
rect 30297 56797 30331 56831
rect 30331 56797 30340 56831
rect 30288 56788 30340 56797
rect 30380 56788 30432 56840
rect 31852 56831 31904 56840
rect 31852 56797 31894 56831
rect 31894 56797 31904 56831
rect 32312 56831 32364 56840
rect 31852 56788 31904 56797
rect 32312 56797 32321 56831
rect 32321 56797 32355 56831
rect 32355 56797 32364 56831
rect 32312 56788 32364 56797
rect 32956 56788 33008 56840
rect 33416 56856 33468 56908
rect 35532 56856 35584 56908
rect 33232 56788 33284 56840
rect 33968 56831 34020 56840
rect 33968 56797 33977 56831
rect 33977 56797 34011 56831
rect 34011 56797 34020 56831
rect 33968 56788 34020 56797
rect 34152 56831 34204 56840
rect 34152 56797 34161 56831
rect 34161 56797 34195 56831
rect 34195 56797 34204 56831
rect 34152 56788 34204 56797
rect 34244 56831 34296 56840
rect 34244 56797 34253 56831
rect 34253 56797 34287 56831
rect 34287 56797 34296 56831
rect 34244 56788 34296 56797
rect 30288 56652 30340 56704
rect 34888 56720 34940 56772
rect 35992 56788 36044 56840
rect 36544 56831 36596 56840
rect 36544 56797 36553 56831
rect 36553 56797 36587 56831
rect 36587 56797 36596 56831
rect 36544 56788 36596 56797
rect 36728 56831 36780 56840
rect 36728 56797 36737 56831
rect 36737 56797 36771 56831
rect 36771 56797 36780 56831
rect 36728 56788 36780 56797
rect 36912 56788 36964 56840
rect 35716 56720 35768 56772
rect 41052 57001 41061 57035
rect 41061 57001 41095 57035
rect 41095 57001 41104 57035
rect 41052 56992 41104 57001
rect 42708 56992 42760 57044
rect 42892 57035 42944 57044
rect 42892 57001 42901 57035
rect 42901 57001 42935 57035
rect 42935 57001 42944 57035
rect 42892 56992 42944 57001
rect 43260 56992 43312 57044
rect 38660 56856 38712 56908
rect 31944 56695 31996 56704
rect 31944 56661 31953 56695
rect 31953 56661 31987 56695
rect 31987 56661 31996 56695
rect 31944 56652 31996 56661
rect 32312 56652 32364 56704
rect 32956 56652 33008 56704
rect 33508 56652 33560 56704
rect 38476 56831 38528 56840
rect 38476 56797 38485 56831
rect 38485 56797 38519 56831
rect 38519 56797 38528 56831
rect 40132 56856 40184 56908
rect 40500 56899 40552 56908
rect 40500 56865 40509 56899
rect 40509 56865 40543 56899
rect 40543 56865 40552 56899
rect 40500 56856 40552 56865
rect 40684 56856 40736 56908
rect 43352 56899 43404 56908
rect 38476 56788 38528 56797
rect 40224 56831 40276 56840
rect 40224 56797 40233 56831
rect 40233 56797 40267 56831
rect 40267 56797 40276 56831
rect 40224 56788 40276 56797
rect 41788 56788 41840 56840
rect 42156 56831 42208 56840
rect 42156 56797 42165 56831
rect 42165 56797 42199 56831
rect 42199 56797 42208 56831
rect 42156 56788 42208 56797
rect 43352 56865 43361 56899
rect 43361 56865 43395 56899
rect 43395 56865 43404 56899
rect 43352 56856 43404 56865
rect 43076 56788 43128 56840
rect 44364 56856 44416 56908
rect 46020 56992 46072 57044
rect 50160 56992 50212 57044
rect 50620 56992 50672 57044
rect 51540 56992 51592 57044
rect 52000 56992 52052 57044
rect 52920 56992 52972 57044
rect 53380 56992 53432 57044
rect 53840 56992 53892 57044
rect 55772 56992 55824 57044
rect 45100 56924 45152 56976
rect 48320 56856 48372 56908
rect 43996 56788 44048 56840
rect 45192 56831 45244 56840
rect 45192 56797 45201 56831
rect 45201 56797 45235 56831
rect 45235 56797 45244 56831
rect 45192 56788 45244 56797
rect 45928 56788 45980 56840
rect 55496 56831 55548 56840
rect 44364 56720 44416 56772
rect 45376 56720 45428 56772
rect 55496 56797 55505 56831
rect 55505 56797 55539 56831
rect 55539 56797 55548 56831
rect 55496 56788 55548 56797
rect 39120 56695 39172 56704
rect 39120 56661 39129 56695
rect 39129 56661 39163 56695
rect 39163 56661 39172 56695
rect 39120 56652 39172 56661
rect 40040 56695 40092 56704
rect 40040 56661 40049 56695
rect 40049 56661 40083 56695
rect 40083 56661 40092 56695
rect 40040 56652 40092 56661
rect 40224 56652 40276 56704
rect 41236 56695 41288 56704
rect 41236 56661 41245 56695
rect 41245 56661 41279 56695
rect 41279 56661 41288 56695
rect 41236 56652 41288 56661
rect 42892 56652 42944 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 23204 56448 23256 56500
rect 23480 56448 23532 56500
rect 26424 56448 26476 56500
rect 27160 56448 27212 56500
rect 27620 56491 27672 56500
rect 27620 56457 27629 56491
rect 27629 56457 27663 56491
rect 27663 56457 27672 56491
rect 27620 56448 27672 56457
rect 27804 56448 27856 56500
rect 29000 56448 29052 56500
rect 30012 56448 30064 56500
rect 30564 56448 30616 56500
rect 30932 56448 30984 56500
rect 31944 56448 31996 56500
rect 32956 56448 33008 56500
rect 34152 56448 34204 56500
rect 35348 56448 35400 56500
rect 38752 56448 38804 56500
rect 5448 56312 5500 56364
rect 22560 56312 22612 56364
rect 23572 56355 23624 56364
rect 23572 56321 23581 56355
rect 23581 56321 23615 56355
rect 23615 56321 23624 56355
rect 23572 56312 23624 56321
rect 23940 56312 23992 56364
rect 25780 56380 25832 56432
rect 25688 56312 25740 56364
rect 28356 56380 28408 56432
rect 27252 56355 27304 56364
rect 23664 56244 23716 56296
rect 25228 56287 25280 56296
rect 25228 56253 25237 56287
rect 25237 56253 25271 56287
rect 25271 56253 25280 56287
rect 25228 56244 25280 56253
rect 17132 56176 17184 56228
rect 26608 56287 26660 56296
rect 26608 56253 26617 56287
rect 26617 56253 26651 56287
rect 26651 56253 26660 56287
rect 26608 56244 26660 56253
rect 27252 56321 27261 56355
rect 27261 56321 27295 56355
rect 27295 56321 27304 56355
rect 27252 56312 27304 56321
rect 27344 56312 27396 56364
rect 28448 56355 28500 56364
rect 27160 56287 27212 56296
rect 27160 56253 27169 56287
rect 27169 56253 27203 56287
rect 27203 56253 27212 56287
rect 27160 56244 27212 56253
rect 28448 56321 28457 56355
rect 28457 56321 28491 56355
rect 28491 56321 28500 56355
rect 28448 56312 28500 56321
rect 29276 56312 29328 56364
rect 29368 56355 29420 56364
rect 29368 56321 29377 56355
rect 29377 56321 29411 56355
rect 29411 56321 29420 56355
rect 29368 56312 29420 56321
rect 29920 56312 29972 56364
rect 31852 56380 31904 56432
rect 33232 56380 33284 56432
rect 32312 56312 32364 56364
rect 32772 56312 32824 56364
rect 32864 56312 32916 56364
rect 30840 56244 30892 56296
rect 31116 56287 31168 56296
rect 31116 56253 31125 56287
rect 31125 56253 31159 56287
rect 31159 56253 31168 56287
rect 33508 56312 33560 56364
rect 34336 56355 34388 56364
rect 34336 56321 34345 56355
rect 34345 56321 34379 56355
rect 34379 56321 34388 56355
rect 34336 56312 34388 56321
rect 35532 56380 35584 56432
rect 36268 56380 36320 56432
rect 36452 56423 36504 56432
rect 36452 56389 36461 56423
rect 36461 56389 36495 56423
rect 36495 56389 36504 56423
rect 36452 56380 36504 56389
rect 36728 56380 36780 56432
rect 37740 56380 37792 56432
rect 42156 56448 42208 56500
rect 42708 56448 42760 56500
rect 43996 56448 44048 56500
rect 39212 56380 39264 56432
rect 39948 56380 40000 56432
rect 40040 56380 40092 56432
rect 35716 56355 35768 56364
rect 35716 56321 35724 56355
rect 35724 56321 35758 56355
rect 35758 56321 35768 56355
rect 35716 56312 35768 56321
rect 35808 56355 35860 56364
rect 35808 56321 35817 56355
rect 35817 56321 35851 56355
rect 35851 56321 35860 56355
rect 35808 56312 35860 56321
rect 36544 56312 36596 56364
rect 36912 56355 36964 56364
rect 36912 56321 36921 56355
rect 36921 56321 36955 56355
rect 36955 56321 36964 56355
rect 36912 56312 36964 56321
rect 31116 56244 31168 56253
rect 34704 56244 34756 56296
rect 38292 56244 38344 56296
rect 39212 56244 39264 56296
rect 31576 56176 31628 56228
rect 34060 56176 34112 56228
rect 34796 56176 34848 56228
rect 34888 56176 34940 56228
rect 35716 56176 35768 56228
rect 39120 56176 39172 56228
rect 40132 56312 40184 56364
rect 40040 56287 40092 56296
rect 40040 56253 40049 56287
rect 40049 56253 40083 56287
rect 40083 56253 40092 56287
rect 40040 56244 40092 56253
rect 40500 56355 40552 56364
rect 40500 56321 40509 56355
rect 40509 56321 40543 56355
rect 40543 56321 40552 56355
rect 40500 56312 40552 56321
rect 40776 56244 40828 56296
rect 42708 56312 42760 56364
rect 43076 56355 43128 56364
rect 41972 56244 42024 56296
rect 42432 56244 42484 56296
rect 42524 56244 42576 56296
rect 43076 56321 43085 56355
rect 43085 56321 43119 56355
rect 43119 56321 43128 56355
rect 43076 56312 43128 56321
rect 43168 56355 43220 56364
rect 43168 56321 43177 56355
rect 43177 56321 43211 56355
rect 43211 56321 43220 56355
rect 43628 56355 43680 56364
rect 43168 56312 43220 56321
rect 43628 56321 43637 56355
rect 43637 56321 43671 56355
rect 43671 56321 43680 56355
rect 43628 56312 43680 56321
rect 43904 56355 43956 56364
rect 43904 56321 43913 56355
rect 43913 56321 43947 56355
rect 43947 56321 43956 56355
rect 45376 56448 45428 56500
rect 49700 56448 49752 56500
rect 51448 56491 51500 56500
rect 51448 56457 51457 56491
rect 51457 56457 51491 56491
rect 51491 56457 51500 56491
rect 51448 56448 51500 56457
rect 53012 56491 53064 56500
rect 53012 56457 53021 56491
rect 53021 56457 53055 56491
rect 53055 56457 53064 56491
rect 53012 56448 53064 56457
rect 54760 56448 54812 56500
rect 55496 56448 55548 56500
rect 43904 56312 43956 56321
rect 43260 56244 43312 56296
rect 45652 56380 45704 56432
rect 44916 56355 44968 56364
rect 44916 56321 44925 56355
rect 44925 56321 44959 56355
rect 44959 56321 44968 56355
rect 44916 56312 44968 56321
rect 45744 56355 45796 56364
rect 45744 56321 45783 56355
rect 45783 56321 45796 56355
rect 45744 56312 45796 56321
rect 44824 56287 44876 56296
rect 44824 56253 44833 56287
rect 44833 56253 44867 56287
rect 44867 56253 44876 56287
rect 44824 56244 44876 56253
rect 46480 56312 46532 56364
rect 47860 56312 47912 56364
rect 48780 56312 48832 56364
rect 49240 56312 49292 56364
rect 46848 56244 46900 56296
rect 39396 56176 39448 56228
rect 44640 56176 44692 56228
rect 25504 56108 25556 56160
rect 25688 56108 25740 56160
rect 32496 56108 32548 56160
rect 33140 56151 33192 56160
rect 33140 56117 33149 56151
rect 33149 56117 33183 56151
rect 33183 56117 33192 56151
rect 33140 56108 33192 56117
rect 33600 56108 33652 56160
rect 34428 56108 34480 56160
rect 35624 56151 35676 56160
rect 35624 56117 35633 56151
rect 35633 56117 35667 56151
rect 35667 56117 35676 56151
rect 35624 56108 35676 56117
rect 36820 56108 36872 56160
rect 37832 56108 37884 56160
rect 40960 56108 41012 56160
rect 41420 56151 41472 56160
rect 41420 56117 41429 56151
rect 41429 56117 41463 56151
rect 41463 56117 41472 56151
rect 41788 56151 41840 56160
rect 41420 56108 41472 56117
rect 41788 56117 41797 56151
rect 41797 56117 41831 56151
rect 41831 56117 41840 56151
rect 41788 56108 41840 56117
rect 43076 56108 43128 56160
rect 45468 56108 45520 56160
rect 45744 56151 45796 56160
rect 45744 56117 45753 56151
rect 45753 56117 45787 56151
rect 45787 56117 45796 56151
rect 45744 56108 45796 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 23756 55904 23808 55956
rect 25044 55904 25096 55956
rect 28448 55904 28500 55956
rect 30380 55904 30432 55956
rect 31576 55947 31628 55956
rect 31576 55913 31585 55947
rect 31585 55913 31619 55947
rect 31619 55913 31628 55947
rect 31576 55904 31628 55913
rect 34428 55904 34480 55956
rect 36912 55904 36964 55956
rect 37832 55904 37884 55956
rect 39120 55904 39172 55956
rect 40132 55904 40184 55956
rect 40500 55904 40552 55956
rect 41880 55904 41932 55956
rect 42708 55904 42760 55956
rect 43168 55904 43220 55956
rect 43444 55947 43496 55956
rect 43444 55913 43453 55947
rect 43453 55913 43487 55947
rect 43487 55913 43496 55947
rect 43444 55904 43496 55913
rect 46848 55947 46900 55956
rect 46848 55913 46857 55947
rect 46857 55913 46891 55947
rect 46891 55913 46900 55947
rect 46848 55904 46900 55913
rect 25228 55768 25280 55820
rect 26516 55768 26568 55820
rect 24032 55743 24084 55752
rect 24032 55709 24041 55743
rect 24041 55709 24075 55743
rect 24075 55709 24084 55743
rect 24032 55700 24084 55709
rect 25596 55700 25648 55752
rect 27344 55700 27396 55752
rect 27160 55564 27212 55616
rect 28356 55700 28408 55752
rect 28448 55632 28500 55684
rect 30012 55768 30064 55820
rect 30748 55768 30800 55820
rect 31116 55768 31168 55820
rect 32496 55836 32548 55888
rect 29000 55700 29052 55752
rect 30932 55743 30984 55752
rect 30932 55709 30941 55743
rect 30941 55709 30975 55743
rect 30975 55709 30984 55743
rect 30932 55700 30984 55709
rect 32772 55768 32824 55820
rect 34704 55836 34756 55888
rect 34888 55879 34940 55888
rect 34888 55845 34897 55879
rect 34897 55845 34931 55879
rect 34931 55845 34940 55879
rect 34888 55836 34940 55845
rect 38200 55836 38252 55888
rect 40960 55836 41012 55888
rect 35164 55811 35216 55820
rect 35164 55777 35173 55811
rect 35173 55777 35207 55811
rect 35207 55777 35216 55811
rect 35164 55768 35216 55777
rect 36820 55811 36872 55820
rect 36820 55777 36829 55811
rect 36829 55777 36863 55811
rect 36863 55777 36872 55811
rect 36820 55768 36872 55777
rect 44364 55879 44416 55888
rect 44364 55845 44373 55879
rect 44373 55845 44407 55879
rect 44407 55845 44416 55879
rect 45468 55879 45520 55888
rect 44364 55836 44416 55845
rect 45468 55845 45477 55879
rect 45477 55845 45511 55879
rect 45511 55845 45520 55879
rect 45468 55836 45520 55845
rect 45652 55836 45704 55888
rect 51816 55768 51868 55820
rect 31392 55743 31444 55752
rect 31392 55709 31401 55743
rect 31401 55709 31435 55743
rect 31435 55709 31444 55743
rect 31392 55700 31444 55709
rect 30104 55675 30156 55684
rect 30104 55641 30113 55675
rect 30113 55641 30147 55675
rect 30147 55641 30156 55675
rect 30104 55632 30156 55641
rect 30288 55675 30340 55684
rect 30288 55641 30297 55675
rect 30297 55641 30331 55675
rect 30331 55641 30340 55675
rect 30288 55632 30340 55641
rect 31024 55632 31076 55684
rect 29276 55564 29328 55616
rect 30012 55564 30064 55616
rect 32588 55700 32640 55752
rect 33140 55743 33192 55752
rect 33140 55709 33149 55743
rect 33149 55709 33183 55743
rect 33183 55709 33192 55743
rect 33140 55700 33192 55709
rect 33232 55700 33284 55752
rect 34060 55743 34112 55752
rect 34060 55709 34069 55743
rect 34069 55709 34103 55743
rect 34103 55709 34112 55743
rect 34060 55700 34112 55709
rect 34244 55700 34296 55752
rect 34428 55700 34480 55752
rect 34612 55700 34664 55752
rect 38200 55700 38252 55752
rect 38568 55743 38620 55752
rect 38568 55709 38577 55743
rect 38577 55709 38611 55743
rect 38611 55709 38620 55743
rect 42524 55743 42576 55752
rect 38568 55700 38620 55709
rect 42524 55709 42533 55743
rect 42533 55709 42567 55743
rect 42567 55709 42576 55743
rect 42524 55700 42576 55709
rect 42892 55700 42944 55752
rect 43996 55700 44048 55752
rect 32404 55675 32456 55684
rect 32404 55641 32413 55675
rect 32413 55641 32447 55675
rect 32447 55641 32456 55675
rect 32404 55632 32456 55641
rect 32864 55632 32916 55684
rect 39396 55675 39448 55684
rect 35348 55564 35400 55616
rect 38476 55607 38528 55616
rect 38476 55573 38485 55607
rect 38485 55573 38519 55607
rect 38519 55573 38528 55607
rect 38476 55564 38528 55573
rect 39396 55641 39405 55675
rect 39405 55641 39439 55675
rect 39439 55641 39448 55675
rect 39396 55632 39448 55641
rect 40224 55675 40276 55684
rect 40224 55641 40233 55675
rect 40233 55641 40267 55675
rect 40267 55641 40276 55675
rect 40224 55632 40276 55641
rect 40408 55675 40460 55684
rect 40408 55641 40417 55675
rect 40417 55641 40451 55675
rect 40451 55641 40460 55675
rect 40408 55632 40460 55641
rect 41880 55632 41932 55684
rect 39304 55564 39356 55616
rect 39488 55564 39540 55616
rect 43628 55632 43680 55684
rect 44824 55700 44876 55752
rect 45376 55743 45428 55752
rect 45376 55709 45385 55743
rect 45385 55709 45419 55743
rect 45419 55709 45428 55743
rect 45376 55700 45428 55709
rect 45744 55632 45796 55684
rect 44916 55564 44968 55616
rect 46204 55607 46256 55616
rect 46204 55573 46213 55607
rect 46213 55573 46247 55607
rect 46247 55573 46256 55607
rect 46204 55564 46256 55573
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 23940 55403 23992 55412
rect 23940 55369 23949 55403
rect 23949 55369 23983 55403
rect 23983 55369 23992 55403
rect 23940 55360 23992 55369
rect 25136 55360 25188 55412
rect 26424 55403 26476 55412
rect 26424 55369 26433 55403
rect 26433 55369 26467 55403
rect 26467 55369 26476 55403
rect 26424 55360 26476 55369
rect 27252 55360 27304 55412
rect 30840 55360 30892 55412
rect 31024 55360 31076 55412
rect 31392 55360 31444 55412
rect 32680 55360 32732 55412
rect 33784 55360 33836 55412
rect 33968 55360 34020 55412
rect 34612 55360 34664 55412
rect 35164 55360 35216 55412
rect 25228 55292 25280 55344
rect 29736 55292 29788 55344
rect 30104 55292 30156 55344
rect 25504 55267 25556 55276
rect 25504 55233 25513 55267
rect 25513 55233 25547 55267
rect 25547 55233 25556 55267
rect 25504 55224 25556 55233
rect 26608 55267 26660 55276
rect 26608 55233 26617 55267
rect 26617 55233 26651 55267
rect 26651 55233 26660 55267
rect 26608 55224 26660 55233
rect 27160 55267 27212 55276
rect 27160 55233 27169 55267
rect 27169 55233 27203 55267
rect 27203 55233 27212 55267
rect 27160 55224 27212 55233
rect 27804 55267 27856 55276
rect 27804 55233 27813 55267
rect 27813 55233 27847 55267
rect 27847 55233 27856 55267
rect 27804 55224 27856 55233
rect 28908 55224 28960 55276
rect 29276 55267 29328 55276
rect 29276 55233 29285 55267
rect 29285 55233 29319 55267
rect 29319 55233 29328 55267
rect 29276 55224 29328 55233
rect 30012 55267 30064 55276
rect 29460 55156 29512 55208
rect 30012 55233 30021 55267
rect 30021 55233 30055 55267
rect 30055 55233 30064 55267
rect 30012 55224 30064 55233
rect 31024 55224 31076 55276
rect 31208 55224 31260 55276
rect 32404 55224 32456 55276
rect 32680 55267 32732 55276
rect 32680 55233 32689 55267
rect 32689 55233 32723 55267
rect 32723 55233 32732 55267
rect 32680 55224 32732 55233
rect 33324 55224 33376 55276
rect 34520 55224 34572 55276
rect 36636 55360 36688 55412
rect 38476 55360 38528 55412
rect 35440 55292 35492 55344
rect 40040 55360 40092 55412
rect 35348 55224 35400 55276
rect 35624 55224 35676 55276
rect 33784 55199 33836 55208
rect 33784 55165 33793 55199
rect 33793 55165 33827 55199
rect 33827 55165 33836 55199
rect 33784 55156 33836 55165
rect 39304 55292 39356 55344
rect 42800 55360 42852 55412
rect 42892 55360 42944 55412
rect 43996 55360 44048 55412
rect 44272 55403 44324 55412
rect 44272 55369 44281 55403
rect 44281 55369 44315 55403
rect 44315 55369 44324 55403
rect 44272 55360 44324 55369
rect 45560 55360 45612 55412
rect 42340 55292 42392 55344
rect 37004 55224 37056 55276
rect 38200 55267 38252 55276
rect 36360 55156 36412 55208
rect 38200 55233 38209 55267
rect 38209 55233 38243 55267
rect 38243 55233 38252 55267
rect 38200 55224 38252 55233
rect 38292 55267 38344 55276
rect 38292 55233 38301 55267
rect 38301 55233 38335 55267
rect 38335 55233 38344 55267
rect 38476 55267 38528 55276
rect 38292 55224 38344 55233
rect 38476 55233 38485 55267
rect 38485 55233 38519 55267
rect 38519 55233 38528 55267
rect 38476 55224 38528 55233
rect 38568 55267 38620 55276
rect 38568 55233 38577 55267
rect 38577 55233 38611 55267
rect 38611 55233 38620 55267
rect 39396 55267 39448 55276
rect 38568 55224 38620 55233
rect 39396 55233 39405 55267
rect 39405 55233 39439 55267
rect 39439 55233 39448 55267
rect 39396 55224 39448 55233
rect 39488 55224 39540 55276
rect 40224 55267 40276 55276
rect 38660 55156 38712 55208
rect 39948 55156 40000 55208
rect 40224 55233 40233 55267
rect 40233 55233 40267 55267
rect 40267 55233 40276 55267
rect 40224 55224 40276 55233
rect 40408 55224 40460 55276
rect 41696 55224 41748 55276
rect 42156 55224 42208 55276
rect 42892 55267 42944 55276
rect 42892 55233 42901 55267
rect 42901 55233 42935 55267
rect 42935 55233 42944 55267
rect 42892 55224 42944 55233
rect 32220 55088 32272 55140
rect 29092 55063 29144 55072
rect 29092 55029 29101 55063
rect 29101 55029 29135 55063
rect 29135 55029 29144 55063
rect 29092 55020 29144 55029
rect 29828 55063 29880 55072
rect 29828 55029 29837 55063
rect 29837 55029 29871 55063
rect 29871 55029 29880 55063
rect 29828 55020 29880 55029
rect 34704 55020 34756 55072
rect 35532 55088 35584 55140
rect 37372 55088 37424 55140
rect 43260 55224 43312 55276
rect 44088 55292 44140 55344
rect 44180 55224 44232 55276
rect 45928 55292 45980 55344
rect 46204 55224 46256 55276
rect 41144 55020 41196 55072
rect 42064 55020 42116 55072
rect 42708 55063 42760 55072
rect 42708 55029 42717 55063
rect 42717 55029 42751 55063
rect 42751 55029 42760 55063
rect 42708 55020 42760 55029
rect 43076 55088 43128 55140
rect 53104 55156 53156 55208
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 25228 54816 25280 54868
rect 25780 54859 25832 54868
rect 25780 54825 25789 54859
rect 25789 54825 25823 54859
rect 25823 54825 25832 54859
rect 25780 54816 25832 54825
rect 26700 54816 26752 54868
rect 28080 54816 28132 54868
rect 29000 54816 29052 54868
rect 30932 54816 30984 54868
rect 31944 54859 31996 54868
rect 31944 54825 31953 54859
rect 31953 54825 31987 54859
rect 31987 54825 31996 54859
rect 31944 54816 31996 54825
rect 32128 54816 32180 54868
rect 33784 54859 33836 54868
rect 33784 54825 33793 54859
rect 33793 54825 33827 54859
rect 33827 54825 33836 54859
rect 33784 54816 33836 54825
rect 34796 54816 34848 54868
rect 35808 54816 35860 54868
rect 37372 54816 37424 54868
rect 38200 54816 38252 54868
rect 40224 54816 40276 54868
rect 40500 54816 40552 54868
rect 41236 54816 41288 54868
rect 41696 54859 41748 54868
rect 41696 54825 41705 54859
rect 41705 54825 41739 54859
rect 41739 54825 41748 54859
rect 41696 54816 41748 54825
rect 28448 54791 28500 54800
rect 28448 54757 28457 54791
rect 28457 54757 28491 54791
rect 28491 54757 28500 54791
rect 28448 54748 28500 54757
rect 35716 54748 35768 54800
rect 36452 54748 36504 54800
rect 37832 54748 37884 54800
rect 40040 54791 40092 54800
rect 40040 54757 40049 54791
rect 40049 54757 40083 54791
rect 40083 54757 40092 54791
rect 40040 54748 40092 54757
rect 25780 54612 25832 54664
rect 27160 54612 27212 54664
rect 29736 54655 29788 54664
rect 29736 54621 29745 54655
rect 29745 54621 29779 54655
rect 29779 54621 29788 54655
rect 29736 54612 29788 54621
rect 29828 54655 29880 54664
rect 29828 54621 29837 54655
rect 29837 54621 29871 54655
rect 29871 54621 29880 54655
rect 29828 54612 29880 54621
rect 28540 54476 28592 54528
rect 29276 54544 29328 54596
rect 30748 54612 30800 54664
rect 31024 54655 31076 54664
rect 31024 54621 31033 54655
rect 31033 54621 31067 54655
rect 31067 54621 31076 54655
rect 31024 54612 31076 54621
rect 31116 54655 31168 54664
rect 31116 54621 31125 54655
rect 31125 54621 31159 54655
rect 31159 54621 31168 54655
rect 31116 54612 31168 54621
rect 31852 54612 31904 54664
rect 32588 54612 32640 54664
rect 33140 54655 33192 54664
rect 33140 54621 33149 54655
rect 33149 54621 33183 54655
rect 33183 54621 33192 54655
rect 33140 54612 33192 54621
rect 39488 54680 39540 54732
rect 41236 54723 41288 54732
rect 41236 54689 41245 54723
rect 41245 54689 41279 54723
rect 41279 54689 41288 54723
rect 42800 54723 42852 54732
rect 41236 54680 41288 54689
rect 39396 54612 39448 54664
rect 33324 54544 33376 54596
rect 33968 54587 34020 54596
rect 33968 54553 33977 54587
rect 33977 54553 34011 54587
rect 34011 54553 34020 54587
rect 33968 54544 34020 54553
rect 34336 54544 34388 54596
rect 42064 54612 42116 54664
rect 42800 54689 42809 54723
rect 42809 54689 42843 54723
rect 42843 54689 42852 54723
rect 42800 54680 42852 54689
rect 43076 54680 43128 54732
rect 43260 54723 43312 54732
rect 43260 54689 43269 54723
rect 43269 54689 43303 54723
rect 43303 54689 43312 54723
rect 43260 54680 43312 54689
rect 44180 54723 44232 54732
rect 44180 54689 44189 54723
rect 44189 54689 44223 54723
rect 44223 54689 44232 54723
rect 44180 54680 44232 54689
rect 43904 54612 43956 54664
rect 29368 54476 29420 54528
rect 32220 54519 32272 54528
rect 32220 54485 32229 54519
rect 32229 54485 32263 54519
rect 32263 54485 32272 54519
rect 32220 54476 32272 54485
rect 32496 54476 32548 54528
rect 42156 54476 42208 54528
rect 42616 54519 42668 54528
rect 42616 54485 42625 54519
rect 42625 54485 42659 54519
rect 42659 54485 42668 54519
rect 42616 54476 42668 54485
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 26516 54315 26568 54324
rect 26516 54281 26525 54315
rect 26525 54281 26559 54315
rect 26559 54281 26568 54315
rect 26516 54272 26568 54281
rect 27160 54315 27212 54324
rect 27160 54281 27169 54315
rect 27169 54281 27203 54315
rect 27203 54281 27212 54315
rect 27160 54272 27212 54281
rect 27804 54315 27856 54324
rect 27804 54281 27813 54315
rect 27813 54281 27847 54315
rect 27847 54281 27856 54315
rect 27804 54272 27856 54281
rect 28264 54315 28316 54324
rect 28264 54281 28273 54315
rect 28273 54281 28307 54315
rect 28307 54281 28316 54315
rect 28264 54272 28316 54281
rect 29276 54272 29328 54324
rect 30748 54272 30800 54324
rect 33232 54272 33284 54324
rect 34336 54315 34388 54324
rect 34336 54281 34345 54315
rect 34345 54281 34379 54315
rect 34379 54281 34388 54315
rect 34336 54272 34388 54281
rect 35532 54272 35584 54324
rect 36452 54315 36504 54324
rect 36452 54281 36461 54315
rect 36461 54281 36495 54315
rect 36495 54281 36504 54315
rect 36452 54272 36504 54281
rect 37280 54272 37332 54324
rect 38936 54272 38988 54324
rect 40500 54315 40552 54324
rect 40500 54281 40509 54315
rect 40509 54281 40543 54315
rect 40543 54281 40552 54315
rect 40500 54272 40552 54281
rect 41788 54272 41840 54324
rect 41972 54315 42024 54324
rect 41972 54281 41981 54315
rect 41981 54281 42015 54315
rect 42015 54281 42024 54315
rect 41972 54272 42024 54281
rect 42708 54315 42760 54324
rect 42708 54281 42717 54315
rect 42717 54281 42751 54315
rect 42751 54281 42760 54315
rect 42708 54272 42760 54281
rect 44180 54315 44232 54324
rect 44180 54281 44189 54315
rect 44189 54281 44223 54315
rect 44223 54281 44232 54315
rect 44180 54272 44232 54281
rect 29092 54136 29144 54188
rect 28540 54111 28592 54120
rect 28540 54077 28549 54111
rect 28549 54077 28583 54111
rect 28583 54077 28592 54111
rect 28540 54068 28592 54077
rect 30288 54136 30340 54188
rect 32680 54204 32732 54256
rect 34520 54204 34572 54256
rect 42156 54204 42208 54256
rect 32496 54179 32548 54188
rect 32496 54145 32505 54179
rect 32505 54145 32539 54179
rect 32539 54145 32548 54179
rect 32496 54136 32548 54145
rect 34060 54136 34112 54188
rect 35348 54136 35400 54188
rect 30104 54068 30156 54120
rect 31024 54068 31076 54120
rect 32220 54068 32272 54120
rect 32588 54068 32640 54120
rect 34152 54068 34204 54120
rect 34704 54068 34756 54120
rect 34796 54068 34848 54120
rect 39580 54136 39632 54188
rect 40316 54179 40368 54188
rect 40316 54145 40325 54179
rect 40325 54145 40359 54179
rect 40359 54145 40368 54179
rect 40316 54136 40368 54145
rect 41144 54179 41196 54188
rect 41144 54145 41153 54179
rect 41153 54145 41187 54179
rect 41187 54145 41196 54179
rect 41144 54136 41196 54145
rect 42616 54179 42668 54188
rect 42616 54145 42625 54179
rect 42625 54145 42659 54179
rect 42659 54145 42668 54179
rect 42616 54136 42668 54145
rect 42984 54136 43036 54188
rect 43260 54136 43312 54188
rect 43996 54179 44048 54188
rect 43996 54145 44005 54179
rect 44005 54145 44039 54179
rect 44039 54145 44048 54179
rect 43996 54136 44048 54145
rect 39948 54068 40000 54120
rect 41236 54111 41288 54120
rect 41236 54077 41245 54111
rect 41245 54077 41279 54111
rect 41279 54077 41288 54111
rect 41236 54068 41288 54077
rect 43076 54068 43128 54120
rect 33324 53932 33376 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 27712 53728 27764 53780
rect 29736 53728 29788 53780
rect 30748 53771 30800 53780
rect 30748 53737 30757 53771
rect 30757 53737 30791 53771
rect 30791 53737 30800 53771
rect 30748 53728 30800 53737
rect 31116 53728 31168 53780
rect 31484 53660 31536 53712
rect 30288 53635 30340 53644
rect 30288 53601 30297 53635
rect 30297 53601 30331 53635
rect 30331 53601 30340 53635
rect 30288 53592 30340 53601
rect 30104 53567 30156 53576
rect 30104 53533 30113 53567
rect 30113 53533 30147 53567
rect 30147 53533 30156 53567
rect 30104 53524 30156 53533
rect 32128 53567 32180 53576
rect 32128 53533 32137 53567
rect 32137 53533 32171 53567
rect 32171 53533 32180 53567
rect 32128 53524 32180 53533
rect 32220 53524 32272 53576
rect 33140 53728 33192 53780
rect 33784 53728 33836 53780
rect 34796 53728 34848 53780
rect 35532 53728 35584 53780
rect 35900 53771 35952 53780
rect 35900 53737 35909 53771
rect 35909 53737 35943 53771
rect 35943 53737 35952 53771
rect 35900 53728 35952 53737
rect 40316 53728 40368 53780
rect 42064 53771 42116 53780
rect 42064 53737 42073 53771
rect 42073 53737 42107 53771
rect 42107 53737 42116 53771
rect 42064 53728 42116 53737
rect 42708 53728 42760 53780
rect 39948 53660 40000 53712
rect 41972 53660 42024 53712
rect 33968 53592 34020 53644
rect 34704 53592 34756 53644
rect 33324 53567 33376 53576
rect 33324 53533 33333 53567
rect 33333 53533 33367 53567
rect 33367 53533 33376 53567
rect 33324 53524 33376 53533
rect 34060 53567 34112 53576
rect 34060 53533 34069 53567
rect 34069 53533 34103 53567
rect 34103 53533 34112 53567
rect 34060 53524 34112 53533
rect 34152 53567 34204 53576
rect 34152 53533 34171 53567
rect 34171 53533 34204 53567
rect 34152 53524 34204 53533
rect 34336 53524 34388 53576
rect 33784 53456 33836 53508
rect 42984 53456 43036 53508
rect 42616 53388 42668 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 30472 53227 30524 53236
rect 30472 53193 30481 53227
rect 30481 53193 30515 53227
rect 30515 53193 30524 53227
rect 30472 53184 30524 53193
rect 31484 53227 31536 53236
rect 31484 53193 31493 53227
rect 31493 53193 31527 53227
rect 31527 53193 31536 53227
rect 31484 53184 31536 53193
rect 32404 53184 32456 53236
rect 39856 53227 39908 53236
rect 39856 53193 39865 53227
rect 39865 53193 39899 53227
rect 39899 53193 39908 53227
rect 39856 53184 39908 53193
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 32036 52640 32088 52692
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 35992 52028 36044 52080
rect 34152 51935 34204 51944
rect 34152 51901 34161 51935
rect 34161 51901 34195 51935
rect 34195 51901 34204 51935
rect 34152 51892 34204 51901
rect 35716 51935 35768 51944
rect 35716 51901 35725 51935
rect 35725 51901 35759 51935
rect 35759 51901 35768 51935
rect 35716 51892 35768 51901
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 34152 51595 34204 51604
rect 34152 51561 34161 51595
rect 34161 51561 34195 51595
rect 34195 51561 34204 51595
rect 34152 51552 34204 51561
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 26516 8576 26568 8628
rect 29000 8576 29052 8628
rect 29828 8576 29880 8628
rect 30104 8236 30156 8288
rect 30656 8304 30708 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 27528 7828 27580 7880
rect 30104 7828 30156 7880
rect 30472 7871 30524 7880
rect 30472 7837 30481 7871
rect 30481 7837 30515 7871
rect 30515 7837 30524 7871
rect 30472 7828 30524 7837
rect 27620 7692 27672 7744
rect 29368 7692 29420 7744
rect 29552 7692 29604 7744
rect 31116 7692 31168 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 29552 7463 29604 7472
rect 29552 7429 29561 7463
rect 29561 7429 29595 7463
rect 29595 7429 29604 7463
rect 29552 7420 29604 7429
rect 30748 7327 30800 7336
rect 30748 7293 30757 7327
rect 30757 7293 30791 7327
rect 30791 7293 30800 7327
rect 30748 7284 30800 7293
rect 27344 7191 27396 7200
rect 27344 7157 27353 7191
rect 27353 7157 27387 7191
rect 27387 7157 27396 7191
rect 27344 7148 27396 7157
rect 27988 7191 28040 7200
rect 27988 7157 27997 7191
rect 27997 7157 28031 7191
rect 28031 7157 28040 7191
rect 27988 7148 28040 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 27344 6851 27396 6860
rect 27344 6817 27353 6851
rect 27353 6817 27387 6851
rect 27387 6817 27396 6851
rect 27344 6808 27396 6817
rect 27620 6808 27672 6860
rect 28080 6851 28132 6860
rect 28080 6817 28089 6851
rect 28089 6817 28123 6851
rect 28123 6817 28132 6851
rect 28080 6808 28132 6817
rect 31116 6851 31168 6860
rect 31116 6817 31125 6851
rect 31125 6817 31159 6851
rect 31159 6817 31168 6851
rect 31116 6808 31168 6817
rect 31668 6851 31720 6860
rect 31668 6817 31677 6851
rect 31677 6817 31711 6851
rect 31711 6817 31720 6851
rect 31668 6808 31720 6817
rect 25228 6604 25280 6656
rect 26424 6740 26476 6792
rect 29828 6740 29880 6792
rect 30932 6783 30984 6792
rect 30932 6749 30941 6783
rect 30941 6749 30975 6783
rect 30975 6749 30984 6783
rect 30932 6740 30984 6749
rect 35348 6740 35400 6792
rect 30104 6672 30156 6724
rect 26516 6604 26568 6656
rect 27344 6604 27396 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 29828 6400 29880 6452
rect 32772 6400 32824 6452
rect 29368 6375 29420 6384
rect 29368 6341 29377 6375
rect 29377 6341 29411 6375
rect 29411 6341 29420 6375
rect 29368 6332 29420 6341
rect 26424 6307 26476 6316
rect 26424 6273 26433 6307
rect 26433 6273 26467 6307
rect 26467 6273 26476 6307
rect 26424 6264 26476 6273
rect 26516 6264 26568 6316
rect 29000 6264 29052 6316
rect 30932 6264 30984 6316
rect 35348 6307 35400 6316
rect 35348 6273 35357 6307
rect 35357 6273 35391 6307
rect 35391 6273 35400 6307
rect 35348 6264 35400 6273
rect 27528 6196 27580 6248
rect 29184 6239 29236 6248
rect 29184 6205 29193 6239
rect 29193 6205 29227 6239
rect 29227 6205 29236 6239
rect 29184 6196 29236 6205
rect 29736 6239 29788 6248
rect 29736 6205 29745 6239
rect 29745 6205 29779 6239
rect 29779 6205 29788 6239
rect 29736 6196 29788 6205
rect 33876 6239 33928 6248
rect 33876 6205 33885 6239
rect 33885 6205 33919 6239
rect 33919 6205 33928 6239
rect 33876 6196 33928 6205
rect 35624 6128 35676 6180
rect 25044 6060 25096 6112
rect 27528 6060 27580 6112
rect 29460 6060 29512 6112
rect 34152 6060 34204 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 35624 5899 35676 5908
rect 35624 5865 35633 5899
rect 35633 5865 35667 5899
rect 35667 5865 35676 5899
rect 35624 5856 35676 5865
rect 25044 5763 25096 5772
rect 25044 5729 25053 5763
rect 25053 5729 25087 5763
rect 25087 5729 25096 5763
rect 25044 5720 25096 5729
rect 25228 5763 25280 5772
rect 25228 5729 25237 5763
rect 25237 5729 25271 5763
rect 25271 5729 25280 5763
rect 25228 5720 25280 5729
rect 25964 5763 26016 5772
rect 25964 5729 25973 5763
rect 25973 5729 26007 5763
rect 26007 5729 26016 5763
rect 25964 5720 26016 5729
rect 27988 5788 28040 5840
rect 27528 5763 27580 5772
rect 27528 5729 27537 5763
rect 27537 5729 27571 5763
rect 27571 5729 27580 5763
rect 27528 5720 27580 5729
rect 27804 5763 27856 5772
rect 27804 5729 27813 5763
rect 27813 5729 27847 5763
rect 27847 5729 27856 5763
rect 27804 5720 27856 5729
rect 30472 5763 30524 5772
rect 30472 5729 30481 5763
rect 30481 5729 30515 5763
rect 30515 5729 30524 5763
rect 30472 5720 30524 5729
rect 30656 5763 30708 5772
rect 30656 5729 30665 5763
rect 30665 5729 30699 5763
rect 30699 5729 30708 5763
rect 30656 5720 30708 5729
rect 31392 5763 31444 5772
rect 31392 5729 31401 5763
rect 31401 5729 31435 5763
rect 31435 5729 31444 5763
rect 31392 5720 31444 5729
rect 29920 5652 29972 5704
rect 32772 5695 32824 5704
rect 32772 5661 32781 5695
rect 32781 5661 32815 5695
rect 32815 5661 32824 5695
rect 32772 5652 32824 5661
rect 35348 5720 35400 5772
rect 34520 5652 34572 5704
rect 33968 5516 34020 5568
rect 36268 5559 36320 5568
rect 36268 5525 36277 5559
rect 36277 5525 36311 5559
rect 36311 5525 36320 5559
rect 36268 5516 36320 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 27344 5287 27396 5296
rect 27344 5253 27353 5287
rect 27353 5253 27387 5287
rect 27387 5253 27396 5287
rect 27344 5244 27396 5253
rect 33968 5287 34020 5296
rect 33968 5253 33977 5287
rect 33977 5253 34011 5287
rect 34011 5253 34020 5287
rect 33968 5244 34020 5253
rect 36268 5287 36320 5296
rect 36268 5253 36277 5287
rect 36277 5253 36311 5287
rect 36311 5253 36320 5287
rect 36268 5244 36320 5253
rect 29460 5219 29512 5228
rect 29460 5185 29469 5219
rect 29469 5185 29503 5219
rect 29503 5185 29512 5219
rect 29460 5176 29512 5185
rect 34152 5219 34204 5228
rect 34152 5185 34161 5219
rect 34161 5185 34195 5219
rect 34195 5185 34204 5219
rect 34152 5176 34204 5185
rect 27712 5151 27764 5160
rect 27712 5117 27721 5151
rect 27721 5117 27755 5151
rect 27755 5117 27764 5151
rect 27712 5108 27764 5117
rect 29644 5151 29696 5160
rect 29644 5117 29653 5151
rect 29653 5117 29687 5151
rect 29687 5117 29696 5151
rect 29644 5108 29696 5117
rect 30380 5151 30432 5160
rect 30380 5117 30389 5151
rect 30389 5117 30423 5151
rect 30423 5117 30432 5151
rect 30380 5108 30432 5117
rect 32496 5151 32548 5160
rect 32496 5117 32505 5151
rect 32505 5117 32539 5151
rect 32539 5117 32548 5151
rect 32496 5108 32548 5117
rect 34704 5151 34756 5160
rect 34704 5117 34713 5151
rect 34713 5117 34747 5151
rect 34747 5117 34756 5151
rect 34704 5108 34756 5117
rect 36452 5151 36504 5160
rect 36452 5117 36461 5151
rect 36461 5117 36495 5151
rect 36495 5117 36504 5151
rect 36452 5108 36504 5117
rect 23664 4972 23716 5024
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 25320 5015 25372 5024
rect 25320 4981 25329 5015
rect 25329 4981 25363 5015
rect 25363 4981 25372 5015
rect 25320 4972 25372 4981
rect 27344 4972 27396 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 23848 4700 23900 4752
rect 21456 4564 21508 4616
rect 22284 4564 22336 4616
rect 23480 4564 23532 4616
rect 26424 4768 26476 4820
rect 29184 4811 29236 4820
rect 29184 4777 29193 4811
rect 29193 4777 29227 4811
rect 29227 4777 29236 4811
rect 29184 4768 29236 4777
rect 36452 4768 36504 4820
rect 26884 4700 26936 4752
rect 25320 4632 25372 4684
rect 27620 4675 27672 4684
rect 27620 4641 27629 4675
rect 27629 4641 27663 4675
rect 27663 4641 27672 4675
rect 27620 4632 27672 4641
rect 29920 4675 29972 4684
rect 29920 4641 29929 4675
rect 29929 4641 29963 4675
rect 29963 4641 29972 4675
rect 29920 4632 29972 4641
rect 30564 4675 30616 4684
rect 30564 4641 30573 4675
rect 30573 4641 30607 4675
rect 30607 4641 30616 4675
rect 30564 4632 30616 4641
rect 32680 4675 32732 4684
rect 32680 4641 32689 4675
rect 32689 4641 32723 4675
rect 32723 4641 32732 4675
rect 32680 4632 32732 4641
rect 34520 4632 34572 4684
rect 26148 4607 26200 4616
rect 26148 4573 26157 4607
rect 26157 4573 26191 4607
rect 26191 4573 26200 4607
rect 26148 4564 26200 4573
rect 35348 4564 35400 4616
rect 35532 4607 35584 4616
rect 35532 4573 35541 4607
rect 35541 4573 35575 4607
rect 35575 4573 35584 4607
rect 35532 4564 35584 4573
rect 36820 4607 36872 4616
rect 36820 4573 36829 4607
rect 36829 4573 36863 4607
rect 36863 4573 36872 4607
rect 36820 4564 36872 4573
rect 30472 4496 30524 4548
rect 26056 4428 26108 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 26148 4224 26200 4276
rect 23480 4131 23532 4140
rect 23480 4097 23489 4131
rect 23489 4097 23523 4131
rect 23523 4097 23532 4131
rect 23480 4088 23532 4097
rect 24676 4088 24728 4140
rect 26884 4088 26936 4140
rect 34612 4088 34664 4140
rect 35348 4088 35400 4140
rect 35624 4088 35676 4140
rect 37372 4088 37424 4140
rect 26424 4063 26476 4072
rect 26424 4029 26433 4063
rect 26433 4029 26467 4063
rect 26467 4029 26476 4063
rect 26424 4020 26476 4029
rect 28356 4063 28408 4072
rect 23112 3952 23164 4004
rect 17316 3884 17368 3936
rect 19432 3884 19484 3936
rect 20352 3884 20404 3936
rect 22008 3884 22060 3936
rect 25320 3952 25372 4004
rect 26056 3952 26108 4004
rect 28356 4029 28365 4063
rect 28365 4029 28399 4063
rect 28399 4029 28408 4063
rect 28356 4020 28408 4029
rect 30840 4063 30892 4072
rect 25872 3884 25924 3936
rect 30840 4029 30849 4063
rect 30849 4029 30883 4063
rect 30883 4029 30892 4063
rect 30840 4020 30892 4029
rect 33048 4063 33100 4072
rect 33048 4029 33057 4063
rect 33057 4029 33091 4063
rect 33091 4029 33100 4063
rect 33048 4020 33100 4029
rect 35532 4020 35584 4072
rect 35808 3952 35860 4004
rect 37188 3952 37240 4004
rect 35440 3884 35492 3936
rect 38292 3884 38344 3936
rect 39396 3884 39448 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 24492 3680 24544 3732
rect 29644 3680 29696 3732
rect 30472 3723 30524 3732
rect 30472 3689 30481 3723
rect 30481 3689 30515 3723
rect 30515 3689 30524 3723
rect 30472 3680 30524 3689
rect 34152 3680 34204 3732
rect 34704 3680 34756 3732
rect 35532 3680 35584 3732
rect 22836 3612 22888 3664
rect 21732 3544 21784 3596
rect 25688 3612 25740 3664
rect 25780 3612 25832 3664
rect 23572 3544 23624 3596
rect 26700 3587 26752 3596
rect 26700 3553 26709 3587
rect 26709 3553 26743 3587
rect 26743 3553 26752 3587
rect 26700 3544 26752 3553
rect 27344 3587 27396 3596
rect 27344 3553 27353 3587
rect 27353 3553 27387 3587
rect 27387 3553 27396 3587
rect 27344 3544 27396 3553
rect 28908 3587 28960 3596
rect 28908 3553 28917 3587
rect 28917 3553 28951 3587
rect 28951 3553 28960 3587
rect 28908 3544 28960 3553
rect 8944 3476 8996 3528
rect 9956 3476 10008 3528
rect 10784 3476 10836 3528
rect 11612 3476 11664 3528
rect 12440 3476 12492 3528
rect 13268 3476 13320 3528
rect 14096 3476 14148 3528
rect 14924 3476 14976 3528
rect 15752 3476 15804 3528
rect 16580 3476 16632 3528
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 18420 3476 18472 3528
rect 19248 3476 19300 3528
rect 20628 3476 20680 3528
rect 23480 3476 23532 3528
rect 23940 3476 23992 3528
rect 30104 3476 30156 3528
rect 34612 3612 34664 3664
rect 36912 3612 36964 3664
rect 39120 3612 39172 3664
rect 41052 3612 41104 3664
rect 45192 3612 45244 3664
rect 47124 3612 47176 3664
rect 32220 3587 32272 3596
rect 32220 3553 32229 3587
rect 32229 3553 32263 3587
rect 32263 3553 32272 3587
rect 32220 3544 32272 3553
rect 33600 3544 33652 3596
rect 36820 3544 36872 3596
rect 39948 3544 40000 3596
rect 41880 3544 41932 3596
rect 42984 3544 43036 3596
rect 37372 3519 37424 3528
rect 37372 3485 37381 3519
rect 37381 3485 37415 3519
rect 37415 3485 37424 3519
rect 37372 3476 37424 3485
rect 24768 3408 24820 3460
rect 30012 3408 30064 3460
rect 30748 3408 30800 3460
rect 34612 3408 34664 3460
rect 37648 3408 37700 3460
rect 40500 3476 40552 3528
rect 42432 3476 42484 3528
rect 44364 3476 44416 3528
rect 45744 3476 45796 3528
rect 46296 3408 46348 3460
rect 47952 3476 48004 3528
rect 49056 3476 49108 3528
rect 50620 3476 50672 3528
rect 50988 3476 51040 3528
rect 51540 3476 51592 3528
rect 36360 3340 36412 3392
rect 40040 3340 40092 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 24032 3136 24084 3188
rect 23940 3068 23992 3120
rect 14372 2932 14424 2984
rect 16304 2932 16356 2984
rect 20904 2932 20956 2984
rect 23296 3000 23348 3052
rect 23756 3000 23808 3052
rect 24032 3000 24084 3052
rect 25780 3136 25832 3188
rect 36912 3136 36964 3188
rect 29000 3068 29052 3120
rect 34796 3068 34848 3120
rect 24308 3000 24360 3052
rect 24584 3000 24636 3052
rect 24768 3043 24820 3052
rect 24768 3009 24777 3043
rect 24777 3009 24811 3043
rect 24811 3009 24820 3043
rect 24768 3000 24820 3009
rect 34704 3000 34756 3052
rect 37372 3000 37424 3052
rect 42708 3000 42760 3052
rect 23480 2932 23532 2984
rect 26976 2932 27028 2984
rect 29184 2975 29236 2984
rect 20076 2864 20128 2916
rect 22560 2864 22612 2916
rect 8208 2796 8260 2848
rect 9680 2796 9732 2848
rect 10232 2796 10284 2848
rect 11060 2796 11112 2848
rect 11336 2796 11388 2848
rect 12716 2796 12768 2848
rect 13544 2796 13596 2848
rect 14648 2796 14700 2848
rect 15476 2796 15528 2848
rect 16856 2796 16908 2848
rect 18144 2796 18196 2848
rect 18696 2796 18748 2848
rect 24584 2796 24636 2848
rect 24860 2796 24912 2848
rect 29184 2941 29193 2975
rect 29193 2941 29227 2975
rect 29227 2941 29236 2975
rect 29184 2932 29236 2941
rect 30104 2975 30156 2984
rect 27896 2864 27948 2916
rect 30104 2941 30113 2975
rect 30113 2941 30147 2975
rect 30147 2941 30156 2975
rect 30104 2932 30156 2941
rect 31116 2975 31168 2984
rect 31116 2941 31125 2975
rect 31125 2941 31159 2975
rect 31159 2941 31168 2975
rect 31116 2932 31168 2941
rect 31944 2932 31996 2984
rect 34428 2932 34480 2984
rect 37464 2932 37516 2984
rect 36084 2864 36136 2916
rect 38844 2932 38896 2984
rect 40776 2932 40828 2984
rect 43260 2932 43312 2984
rect 37740 2864 37792 2916
rect 29460 2796 29512 2848
rect 30196 2796 30248 2848
rect 37556 2839 37608 2848
rect 37556 2805 37565 2839
rect 37565 2805 37599 2839
rect 37599 2805 37608 2839
rect 37556 2796 37608 2805
rect 39672 2864 39724 2916
rect 41604 2864 41656 2916
rect 44916 2864 44968 2916
rect 48780 2932 48832 2984
rect 43812 2796 43864 2848
rect 45468 2796 45520 2848
rect 47676 2864 47728 2916
rect 49608 2864 49660 2916
rect 50712 2864 50764 2916
rect 46848 2796 46900 2848
rect 48228 2796 48280 2848
rect 50160 2796 50212 2848
rect 52092 2796 52144 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 23480 2592 23532 2644
rect 24860 2592 24912 2644
rect 8576 2524 8628 2576
rect 10508 2524 10560 2576
rect 15200 2524 15252 2576
rect 17132 2524 17184 2576
rect 18972 2524 19024 2576
rect 23572 2524 23624 2576
rect 13820 2456 13872 2508
rect 17868 2456 17920 2508
rect 19984 2456 20036 2508
rect 23388 2456 23440 2508
rect 24584 2456 24636 2508
rect 7656 2388 7708 2440
rect 9312 2388 9364 2440
rect 12164 2388 12216 2440
rect 12992 2388 13044 2440
rect 16028 2388 16080 2440
rect 11888 2320 11940 2372
rect 21180 2320 21232 2372
rect 23296 2388 23348 2440
rect 24032 2431 24084 2440
rect 24032 2397 24041 2431
rect 24041 2397 24075 2431
rect 24075 2397 24084 2431
rect 24032 2388 24084 2397
rect 25780 2431 25832 2440
rect 25780 2397 25789 2431
rect 25789 2397 25823 2431
rect 25823 2397 25832 2431
rect 25780 2388 25832 2397
rect 25872 2388 25924 2440
rect 28540 2499 28592 2508
rect 28540 2465 28549 2499
rect 28549 2465 28583 2499
rect 28583 2465 28592 2499
rect 28540 2456 28592 2465
rect 34612 2592 34664 2644
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 38752 2635 38804 2644
rect 38752 2601 38761 2635
rect 38761 2601 38795 2635
rect 38795 2601 38804 2635
rect 38752 2592 38804 2601
rect 40040 2635 40092 2644
rect 40040 2601 40049 2635
rect 40049 2601 40083 2635
rect 40083 2601 40092 2635
rect 40040 2592 40092 2601
rect 34704 2524 34756 2576
rect 42156 2524 42208 2576
rect 44640 2524 44692 2576
rect 48504 2524 48556 2576
rect 51816 2524 51868 2576
rect 30196 2499 30248 2508
rect 30196 2465 30205 2499
rect 30205 2465 30239 2499
rect 30239 2465 30248 2499
rect 30196 2456 30248 2465
rect 33324 2499 33376 2508
rect 33324 2465 33333 2499
rect 33333 2465 33367 2499
rect 33367 2465 33376 2499
rect 33324 2456 33376 2465
rect 35440 2456 35492 2508
rect 38016 2456 38068 2508
rect 41420 2456 41472 2508
rect 43536 2456 43588 2508
rect 46572 2456 46624 2508
rect 49332 2456 49384 2508
rect 52368 2456 52420 2508
rect 25596 2320 25648 2372
rect 35624 2388 35676 2440
rect 27896 2320 27948 2372
rect 29000 2320 29052 2372
rect 34704 2320 34756 2372
rect 34796 2320 34848 2372
rect 25044 2252 25096 2304
rect 30104 2252 30156 2304
rect 34980 2252 35032 2304
rect 38568 2388 38620 2440
rect 40224 2320 40276 2372
rect 44088 2320 44140 2372
rect 46020 2388 46072 2440
rect 47400 2320 47452 2372
rect 49884 2388 49936 2440
rect 51264 2320 51316 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 34704 2048 34756 2100
rect 37556 2048 37608 2100
rect 23756 1436 23808 1488
rect 24216 1436 24268 1488
rect 34704 1368 34756 1420
rect 35716 1368 35768 1420
<< metal2 >>
rect 3698 59200 3754 60000
rect 4158 59200 4214 60000
rect 4618 59200 4674 60000
rect 5078 59200 5134 60000
rect 5538 59200 5594 60000
rect 5998 59200 6054 60000
rect 6458 59200 6514 60000
rect 6918 59200 6974 60000
rect 7378 59200 7434 60000
rect 7838 59200 7894 60000
rect 8298 59200 8354 60000
rect 8758 59200 8814 60000
rect 9218 59200 9274 60000
rect 9678 59200 9734 60000
rect 10138 59200 10194 60000
rect 10598 59200 10654 60000
rect 11058 59200 11114 60000
rect 11518 59200 11574 60000
rect 11978 59200 12034 60000
rect 12438 59200 12494 60000
rect 12898 59200 12954 60000
rect 13358 59200 13414 60000
rect 13818 59200 13874 60000
rect 14278 59200 14334 60000
rect 14738 59200 14794 60000
rect 15198 59200 15254 60000
rect 15658 59200 15714 60000
rect 16118 59200 16174 60000
rect 16578 59200 16634 60000
rect 17038 59200 17094 60000
rect 17498 59200 17554 60000
rect 17958 59200 18014 60000
rect 18418 59200 18474 60000
rect 18878 59200 18934 60000
rect 18984 59214 19288 59242
rect 3712 57594 3740 59200
rect 3700 57588 3752 57594
rect 3700 57530 3752 57536
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4632 57050 4660 59200
rect 5092 57594 5120 59200
rect 5080 57588 5132 57594
rect 5080 57530 5132 57536
rect 5448 57316 5500 57322
rect 5448 57258 5500 57264
rect 4620 57044 4672 57050
rect 4620 56986 4672 56992
rect 5460 56370 5488 57258
rect 6012 57050 6040 59200
rect 6092 57384 6144 57390
rect 6090 57352 6092 57361
rect 6144 57352 6146 57361
rect 6090 57287 6146 57296
rect 6472 57050 6500 59200
rect 7392 57458 7420 59200
rect 7852 57458 7880 59200
rect 8772 57458 8800 59200
rect 9232 57458 9260 59200
rect 10152 57458 10180 59200
rect 10612 57594 10640 59200
rect 10600 57588 10652 57594
rect 10600 57530 10652 57536
rect 7380 57452 7432 57458
rect 7380 57394 7432 57400
rect 7840 57452 7892 57458
rect 7840 57394 7892 57400
rect 8760 57452 8812 57458
rect 8760 57394 8812 57400
rect 9220 57452 9272 57458
rect 9220 57394 9272 57400
rect 10140 57452 10192 57458
rect 10140 57394 10192 57400
rect 10968 57452 11020 57458
rect 10968 57394 11020 57400
rect 6000 57044 6052 57050
rect 6000 56986 6052 56992
rect 6460 57044 6512 57050
rect 6460 56986 6512 56992
rect 10980 56982 11008 57394
rect 11532 57050 11560 59200
rect 11992 57594 12020 59200
rect 11980 57588 12032 57594
rect 11980 57530 12032 57536
rect 12346 57488 12402 57497
rect 12912 57458 12940 59200
rect 13372 57594 13400 59200
rect 13360 57588 13412 57594
rect 13360 57530 13412 57536
rect 12346 57423 12348 57432
rect 12400 57423 12402 57432
rect 12900 57452 12952 57458
rect 12348 57394 12400 57400
rect 12900 57394 12952 57400
rect 14292 57050 14320 59200
rect 14752 57594 14780 59200
rect 14740 57588 14792 57594
rect 14740 57530 14792 57536
rect 15672 57458 15700 59200
rect 16132 57594 16160 59200
rect 16120 57588 16172 57594
rect 16120 57530 16172 57536
rect 15660 57452 15712 57458
rect 15660 57394 15712 57400
rect 17052 57050 17080 59200
rect 17512 57594 17540 59200
rect 17868 57860 17920 57866
rect 17868 57802 17920 57808
rect 17500 57588 17552 57594
rect 17500 57530 17552 57536
rect 17880 57458 17908 57802
rect 18432 57458 18460 59200
rect 18892 59106 18920 59200
rect 18984 59106 19012 59214
rect 18892 59078 19012 59106
rect 19260 57610 19288 59214
rect 19338 59200 19394 60000
rect 19798 59200 19854 60000
rect 20258 59200 20314 60000
rect 20718 59200 20774 60000
rect 21178 59200 21234 60000
rect 21638 59200 21694 60000
rect 22098 59200 22154 60000
rect 22558 59200 22614 60000
rect 23018 59200 23074 60000
rect 23478 59200 23534 60000
rect 23938 59200 23994 60000
rect 24398 59200 24454 60000
rect 24858 59200 24914 60000
rect 25318 59200 25374 60000
rect 25778 59200 25834 60000
rect 26238 59200 26294 60000
rect 26698 59200 26754 60000
rect 27158 59200 27214 60000
rect 27618 59200 27674 60000
rect 28078 59200 28134 60000
rect 28538 59200 28594 60000
rect 28998 59200 29054 60000
rect 29458 59200 29514 60000
rect 29918 59200 29974 60000
rect 30378 59200 30434 60000
rect 30838 59200 30894 60000
rect 31298 59200 31354 60000
rect 31758 59200 31814 60000
rect 31864 59214 32076 59242
rect 19812 58018 19840 59200
rect 19812 57990 20024 58018
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 19260 57594 19380 57610
rect 19260 57588 19392 57594
rect 19260 57582 19340 57588
rect 19340 57530 19392 57536
rect 17132 57452 17184 57458
rect 17132 57394 17184 57400
rect 17868 57452 17920 57458
rect 17868 57394 17920 57400
rect 18420 57452 18472 57458
rect 18420 57394 18472 57400
rect 11520 57044 11572 57050
rect 11520 56986 11572 56992
rect 14280 57044 14332 57050
rect 14280 56986 14332 56992
rect 17040 57044 17092 57050
rect 17040 56986 17092 56992
rect 10968 56976 11020 56982
rect 10968 56918 11020 56924
rect 5448 56364 5500 56370
rect 5448 56306 5500 56312
rect 17144 56234 17172 57394
rect 19996 57050 20024 57990
rect 20272 57594 20300 59200
rect 20260 57588 20312 57594
rect 20260 57530 20312 57536
rect 21192 57050 21220 59200
rect 21364 57928 21416 57934
rect 21364 57870 21416 57876
rect 19984 57044 20036 57050
rect 19984 56986 20036 56992
rect 21180 57044 21232 57050
rect 21180 56986 21232 56992
rect 21376 56982 21404 57870
rect 21652 57050 21680 59200
rect 22192 57588 22244 57594
rect 22192 57530 22244 57536
rect 21640 57044 21692 57050
rect 21640 56986 21692 56992
rect 21364 56976 21416 56982
rect 21364 56918 21416 56924
rect 22204 56778 22232 57530
rect 22192 56772 22244 56778
rect 22192 56714 22244 56720
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 22572 56370 22600 59200
rect 22836 57792 22888 57798
rect 22836 57734 22888 57740
rect 22744 57384 22796 57390
rect 22744 57326 22796 57332
rect 22756 56914 22784 57326
rect 22848 57254 22876 57734
rect 23032 57594 23060 59200
rect 23952 57798 23980 59200
rect 23940 57792 23992 57798
rect 23940 57734 23992 57740
rect 23020 57588 23072 57594
rect 23020 57530 23072 57536
rect 24412 57526 24440 59200
rect 24768 57792 24820 57798
rect 24768 57734 24820 57740
rect 23480 57520 23532 57526
rect 23480 57462 23532 57468
rect 24400 57520 24452 57526
rect 24400 57462 24452 57468
rect 23204 57452 23256 57458
rect 23204 57394 23256 57400
rect 22836 57248 22888 57254
rect 22836 57190 22888 57196
rect 23216 57050 23244 57394
rect 23492 57322 23520 57462
rect 24780 57458 24808 57734
rect 25044 57588 25096 57594
rect 25044 57530 25096 57536
rect 23664 57452 23716 57458
rect 23664 57394 23716 57400
rect 23756 57452 23808 57458
rect 23756 57394 23808 57400
rect 24768 57452 24820 57458
rect 24768 57394 24820 57400
rect 23480 57316 23532 57322
rect 23480 57258 23532 57264
rect 23572 57316 23624 57322
rect 23572 57258 23624 57264
rect 23204 57044 23256 57050
rect 23204 56986 23256 56992
rect 22744 56908 22796 56914
rect 22744 56850 22796 56856
rect 23216 56506 23244 56986
rect 23480 56840 23532 56846
rect 23480 56782 23532 56788
rect 23492 56506 23520 56782
rect 23204 56500 23256 56506
rect 23204 56442 23256 56448
rect 23480 56500 23532 56506
rect 23480 56442 23532 56448
rect 23584 56370 23612 57258
rect 22560 56364 22612 56370
rect 22560 56306 22612 56312
rect 23572 56364 23624 56370
rect 23572 56306 23624 56312
rect 23676 56302 23704 57394
rect 23768 57338 23796 57394
rect 23768 57310 23980 57338
rect 23848 57248 23900 57254
rect 23848 57190 23900 57196
rect 23860 57050 23888 57190
rect 23848 57044 23900 57050
rect 23848 56986 23900 56992
rect 23756 56908 23808 56914
rect 23756 56850 23808 56856
rect 23664 56296 23716 56302
rect 23664 56238 23716 56244
rect 17132 56228 17184 56234
rect 17132 56170 17184 56176
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 23768 55962 23796 56850
rect 23846 56808 23902 56817
rect 23952 56794 23980 57310
rect 24032 57248 24084 57254
rect 24032 57190 24084 57196
rect 24124 57248 24176 57254
rect 24124 57190 24176 57196
rect 23902 56766 23980 56794
rect 23846 56743 23902 56752
rect 23860 56710 23888 56743
rect 23848 56704 23900 56710
rect 23848 56646 23900 56652
rect 23940 56364 23992 56370
rect 23940 56306 23992 56312
rect 23756 55956 23808 55962
rect 23756 55898 23808 55904
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 23952 55418 23980 56306
rect 24044 55758 24072 57190
rect 24136 56982 24164 57190
rect 24124 56976 24176 56982
rect 24124 56918 24176 56924
rect 24780 56846 24808 57394
rect 25056 56914 25084 57530
rect 25136 57452 25188 57458
rect 25136 57394 25188 57400
rect 25044 56908 25096 56914
rect 25044 56850 25096 56856
rect 24768 56840 24820 56846
rect 24768 56782 24820 56788
rect 25056 55962 25084 56850
rect 25148 56846 25176 57394
rect 25228 57384 25280 57390
rect 25228 57326 25280 57332
rect 25136 56840 25188 56846
rect 25136 56782 25188 56788
rect 25044 55956 25096 55962
rect 25044 55898 25096 55904
rect 24032 55752 24084 55758
rect 24032 55694 24084 55700
rect 25148 55418 25176 56782
rect 25240 56302 25268 57326
rect 25332 57254 25360 59200
rect 25792 57594 25820 59200
rect 25780 57588 25832 57594
rect 25780 57530 25832 57536
rect 25320 57248 25372 57254
rect 25320 57190 25372 57196
rect 25688 56840 25740 56846
rect 25688 56782 25740 56788
rect 25596 56704 25648 56710
rect 25596 56646 25648 56652
rect 25228 56296 25280 56302
rect 25228 56238 25280 56244
rect 25240 55826 25268 56238
rect 25504 56160 25556 56166
rect 25504 56102 25556 56108
rect 25228 55820 25280 55826
rect 25228 55762 25280 55768
rect 23940 55412 23992 55418
rect 23940 55354 23992 55360
rect 25136 55412 25188 55418
rect 25136 55354 25188 55360
rect 25240 55350 25268 55762
rect 25228 55344 25280 55350
rect 25228 55286 25280 55292
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 25240 54874 25268 55286
rect 25516 55282 25544 56102
rect 25608 55865 25636 56646
rect 25700 56370 25728 56782
rect 26424 56500 26476 56506
rect 26424 56442 26476 56448
rect 25780 56432 25832 56438
rect 25780 56374 25832 56380
rect 25688 56364 25740 56370
rect 25688 56306 25740 56312
rect 25700 56166 25728 56306
rect 25688 56160 25740 56166
rect 25688 56102 25740 56108
rect 25594 55856 25650 55865
rect 25594 55791 25650 55800
rect 25608 55758 25636 55791
rect 25596 55752 25648 55758
rect 25596 55694 25648 55700
rect 25504 55276 25556 55282
rect 25504 55218 25556 55224
rect 25792 54874 25820 56374
rect 26436 55418 26464 56442
rect 26608 56296 26660 56302
rect 26608 56238 26660 56244
rect 26516 55820 26568 55826
rect 26516 55762 26568 55768
rect 26424 55412 26476 55418
rect 26424 55354 26476 55360
rect 25228 54868 25280 54874
rect 25228 54810 25280 54816
rect 25780 54868 25832 54874
rect 25780 54810 25832 54816
rect 25792 54670 25820 54810
rect 25780 54664 25832 54670
rect 25780 54606 25832 54612
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 26528 54330 26556 55762
rect 26620 55282 26648 56238
rect 26608 55276 26660 55282
rect 26608 55218 26660 55224
rect 26712 54874 26740 59200
rect 27172 57594 27200 59200
rect 27436 57928 27488 57934
rect 27436 57870 27488 57876
rect 27160 57588 27212 57594
rect 27160 57530 27212 57536
rect 27252 57452 27304 57458
rect 27252 57394 27304 57400
rect 27158 57352 27214 57361
rect 27158 57287 27214 57296
rect 27172 57050 27200 57287
rect 27160 57044 27212 57050
rect 27160 56986 27212 56992
rect 27160 56500 27212 56506
rect 27160 56442 27212 56448
rect 27172 56302 27200 56442
rect 27264 56370 27292 57394
rect 27448 57050 27476 57870
rect 27526 57488 27582 57497
rect 27526 57423 27582 57432
rect 27436 57044 27488 57050
rect 27436 56986 27488 56992
rect 27448 56846 27476 56986
rect 27540 56846 27568 57423
rect 27620 57044 27672 57050
rect 27672 57004 27752 57032
rect 27620 56986 27672 56992
rect 27436 56840 27488 56846
rect 27436 56782 27488 56788
rect 27528 56840 27580 56846
rect 27528 56782 27580 56788
rect 27540 56710 27568 56782
rect 27528 56704 27580 56710
rect 27528 56646 27580 56652
rect 27620 56500 27672 56506
rect 27620 56442 27672 56448
rect 27252 56364 27304 56370
rect 27252 56306 27304 56312
rect 27344 56364 27396 56370
rect 27344 56306 27396 56312
rect 27160 56296 27212 56302
rect 27160 56238 27212 56244
rect 27160 55616 27212 55622
rect 27160 55558 27212 55564
rect 27172 55282 27200 55558
rect 27264 55418 27292 56306
rect 27356 55758 27384 56306
rect 27632 56273 27660 56442
rect 27618 56264 27674 56273
rect 27618 56199 27674 56208
rect 27344 55752 27396 55758
rect 27344 55694 27396 55700
rect 27252 55412 27304 55418
rect 27252 55354 27304 55360
rect 27160 55276 27212 55282
rect 27160 55218 27212 55224
rect 26700 54868 26752 54874
rect 26700 54810 26752 54816
rect 27160 54664 27212 54670
rect 27160 54606 27212 54612
rect 27172 54330 27200 54606
rect 26516 54324 26568 54330
rect 26516 54266 26568 54272
rect 27160 54324 27212 54330
rect 27160 54266 27212 54272
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 26528 8634 26556 54266
rect 27724 53786 27752 57004
rect 27804 56840 27856 56846
rect 27804 56782 27856 56788
rect 27816 56506 27844 56782
rect 27804 56500 27856 56506
rect 27804 56442 27856 56448
rect 27804 55276 27856 55282
rect 27804 55218 27856 55224
rect 27816 54330 27844 55218
rect 28092 54874 28120 59200
rect 28448 57860 28500 57866
rect 28448 57802 28500 57808
rect 28460 56982 28488 57802
rect 28552 57594 28580 59200
rect 29012 57610 29040 59200
rect 29184 57792 29236 57798
rect 29184 57734 29236 57740
rect 28540 57588 28592 57594
rect 29012 57582 29132 57610
rect 28540 57530 28592 57536
rect 28816 57248 28868 57254
rect 28816 57190 28868 57196
rect 28908 57248 28960 57254
rect 28908 57190 28960 57196
rect 28828 56982 28856 57190
rect 28920 57050 28948 57190
rect 28908 57044 28960 57050
rect 28908 56986 28960 56992
rect 28356 56976 28408 56982
rect 28356 56918 28408 56924
rect 28448 56976 28500 56982
rect 28448 56918 28500 56924
rect 28816 56976 28868 56982
rect 28816 56918 28868 56924
rect 28264 56908 28316 56914
rect 28264 56850 28316 56856
rect 28080 54868 28132 54874
rect 28080 54810 28132 54816
rect 28276 54330 28304 56850
rect 28368 56438 28396 56918
rect 28724 56704 28776 56710
rect 28776 56664 29040 56692
rect 28724 56646 28776 56652
rect 29012 56506 29040 56664
rect 29000 56500 29052 56506
rect 29000 56442 29052 56448
rect 28356 56432 28408 56438
rect 28356 56374 28408 56380
rect 28368 55758 28396 56374
rect 28448 56364 28500 56370
rect 28448 56306 28500 56312
rect 28460 55962 28488 56306
rect 28448 55956 28500 55962
rect 28448 55898 28500 55904
rect 29104 55842 29132 57582
rect 29196 57526 29224 57734
rect 29184 57520 29236 57526
rect 29184 57462 29236 57468
rect 29196 56846 29224 57462
rect 29276 57452 29328 57458
rect 29276 57394 29328 57400
rect 29288 56914 29316 57394
rect 29276 56908 29328 56914
rect 29276 56850 29328 56856
rect 29184 56840 29236 56846
rect 29184 56782 29236 56788
rect 29366 56400 29422 56409
rect 29276 56364 29328 56370
rect 29366 56335 29368 56344
rect 29276 56306 29328 56312
rect 29420 56335 29422 56344
rect 29368 56306 29420 56312
rect 28920 55814 29132 55842
rect 28356 55752 28408 55758
rect 28356 55694 28408 55700
rect 28448 55684 28500 55690
rect 28448 55626 28500 55632
rect 28460 54806 28488 55626
rect 28920 55282 28948 55814
rect 29000 55752 29052 55758
rect 29000 55694 29052 55700
rect 28908 55276 28960 55282
rect 28908 55218 28960 55224
rect 29012 54874 29040 55694
rect 29288 55622 29316 56306
rect 29276 55616 29328 55622
rect 29276 55558 29328 55564
rect 29276 55276 29328 55282
rect 29276 55218 29328 55224
rect 29092 55072 29144 55078
rect 29092 55014 29144 55020
rect 29000 54868 29052 54874
rect 29000 54810 29052 54816
rect 28448 54800 28500 54806
rect 28448 54742 28500 54748
rect 28540 54528 28592 54534
rect 28540 54470 28592 54476
rect 27804 54324 27856 54330
rect 27804 54266 27856 54272
rect 28264 54324 28316 54330
rect 28264 54266 28316 54272
rect 28552 54126 28580 54470
rect 29104 54194 29132 55014
rect 29288 54602 29316 55218
rect 29276 54596 29328 54602
rect 29276 54538 29328 54544
rect 29288 54330 29316 54538
rect 29380 54534 29408 56306
rect 29472 55214 29500 59200
rect 29932 56370 29960 59200
rect 30392 57474 30420 59200
rect 30564 57860 30616 57866
rect 30564 57802 30616 57808
rect 30392 57458 30512 57474
rect 30392 57452 30524 57458
rect 30392 57446 30472 57452
rect 30472 57394 30524 57400
rect 30012 57384 30064 57390
rect 30012 57326 30064 57332
rect 30024 56914 30052 57326
rect 30288 57316 30340 57322
rect 30288 57258 30340 57264
rect 30012 56908 30064 56914
rect 30012 56850 30064 56856
rect 30300 56846 30328 57258
rect 30288 56840 30340 56846
rect 30288 56782 30340 56788
rect 30380 56840 30432 56846
rect 30380 56782 30432 56788
rect 30012 56772 30064 56778
rect 30012 56714 30064 56720
rect 30024 56506 30052 56714
rect 30300 56710 30328 56782
rect 30288 56704 30340 56710
rect 30288 56646 30340 56652
rect 30012 56500 30064 56506
rect 30012 56442 30064 56448
rect 29920 56364 29972 56370
rect 29920 56306 29972 56312
rect 30024 55826 30052 56442
rect 30392 55962 30420 56782
rect 30380 55956 30432 55962
rect 30380 55898 30432 55904
rect 30012 55820 30064 55826
rect 30012 55762 30064 55768
rect 30286 55720 30342 55729
rect 30104 55684 30156 55690
rect 30286 55655 30288 55664
rect 30104 55626 30156 55632
rect 30340 55655 30342 55664
rect 30288 55626 30340 55632
rect 30012 55616 30064 55622
rect 30012 55558 30064 55564
rect 29736 55344 29788 55350
rect 29736 55286 29788 55292
rect 29460 55208 29512 55214
rect 29460 55150 29512 55156
rect 29748 54670 29776 55286
rect 30024 55282 30052 55558
rect 30116 55350 30144 55626
rect 30104 55344 30156 55350
rect 30104 55286 30156 55292
rect 30012 55276 30064 55282
rect 30012 55218 30064 55224
rect 29828 55072 29880 55078
rect 29828 55014 29880 55020
rect 29840 54670 29868 55014
rect 29736 54664 29788 54670
rect 29736 54606 29788 54612
rect 29828 54664 29880 54670
rect 29828 54606 29880 54612
rect 29368 54528 29420 54534
rect 29368 54470 29420 54476
rect 29276 54324 29328 54330
rect 29276 54266 29328 54272
rect 29092 54188 29144 54194
rect 29092 54130 29144 54136
rect 28540 54120 28592 54126
rect 28540 54062 28592 54068
rect 29748 53786 29776 54606
rect 30288 54188 30340 54194
rect 30288 54130 30340 54136
rect 30104 54120 30156 54126
rect 30104 54062 30156 54068
rect 27712 53780 27764 53786
rect 27712 53722 27764 53728
rect 29736 53780 29788 53786
rect 29736 53722 29788 53728
rect 30116 53582 30144 54062
rect 30300 53650 30328 54130
rect 30288 53644 30340 53650
rect 30288 53586 30340 53592
rect 30104 53576 30156 53582
rect 30104 53518 30156 53524
rect 30484 53242 30512 57394
rect 30576 56506 30604 57802
rect 30852 57458 30880 59200
rect 30840 57452 30892 57458
rect 30840 57394 30892 57400
rect 31312 57050 31340 59200
rect 31772 59106 31800 59200
rect 31864 59106 31892 59214
rect 31772 59078 31892 59106
rect 31576 57520 31628 57526
rect 31576 57462 31628 57468
rect 31588 57254 31616 57462
rect 32048 57390 32076 59214
rect 32218 59200 32274 60000
rect 32678 59200 32734 60000
rect 33138 59200 33194 60000
rect 33598 59200 33654 60000
rect 34058 59200 34114 60000
rect 34518 59200 34574 60000
rect 34978 59200 35034 60000
rect 35084 59214 35388 59242
rect 31852 57384 31904 57390
rect 31852 57326 31904 57332
rect 32036 57384 32088 57390
rect 32036 57326 32088 57332
rect 31576 57248 31628 57254
rect 31576 57190 31628 57196
rect 31300 57044 31352 57050
rect 31300 56986 31352 56992
rect 31864 56846 31892 57326
rect 31944 56976 31996 56982
rect 31944 56918 31996 56924
rect 31852 56840 31904 56846
rect 31852 56782 31904 56788
rect 30564 56500 30616 56506
rect 30932 56500 30984 56506
rect 30564 56442 30616 56448
rect 30852 56460 30932 56488
rect 30852 56302 30880 56460
rect 30932 56442 30984 56448
rect 31864 56438 31892 56782
rect 31956 56710 31984 56918
rect 31944 56704 31996 56710
rect 31944 56646 31996 56652
rect 31956 56506 31984 56646
rect 31944 56500 31996 56506
rect 31944 56442 31996 56448
rect 31852 56432 31904 56438
rect 31852 56374 31904 56380
rect 30840 56296 30892 56302
rect 30840 56238 30892 56244
rect 31116 56296 31168 56302
rect 31116 56238 31168 56244
rect 30748 55820 30800 55826
rect 30748 55762 30800 55768
rect 30760 54670 30788 55762
rect 30852 55418 30880 56238
rect 31128 55826 31156 56238
rect 31576 56228 31628 56234
rect 31576 56170 31628 56176
rect 31588 55962 31616 56170
rect 31576 55956 31628 55962
rect 31576 55898 31628 55904
rect 31116 55820 31168 55826
rect 31116 55762 31168 55768
rect 30932 55752 30984 55758
rect 30932 55694 30984 55700
rect 31392 55752 31444 55758
rect 31392 55694 31444 55700
rect 30840 55412 30892 55418
rect 30840 55354 30892 55360
rect 30944 54874 30972 55694
rect 31024 55684 31076 55690
rect 31024 55626 31076 55632
rect 31036 55418 31064 55626
rect 31404 55418 31432 55694
rect 31024 55412 31076 55418
rect 31024 55354 31076 55360
rect 31392 55412 31444 55418
rect 31392 55354 31444 55360
rect 31024 55276 31076 55282
rect 31024 55218 31076 55224
rect 31208 55276 31260 55282
rect 31208 55218 31260 55224
rect 30932 54868 30984 54874
rect 30932 54810 30984 54816
rect 31036 54670 31064 55218
rect 30748 54664 30800 54670
rect 30748 54606 30800 54612
rect 31024 54664 31076 54670
rect 31024 54606 31076 54612
rect 31116 54664 31168 54670
rect 31220 54652 31248 55218
rect 31864 54670 31892 56374
rect 31956 54874 31984 56442
rect 31944 54868 31996 54874
rect 31944 54810 31996 54816
rect 31168 54624 31248 54652
rect 31852 54664 31904 54670
rect 31116 54606 31168 54612
rect 31852 54606 31904 54612
rect 30760 54330 30788 54606
rect 30748 54324 30800 54330
rect 30748 54266 30800 54272
rect 30760 53786 30788 54266
rect 31036 54126 31064 54606
rect 31024 54120 31076 54126
rect 31024 54062 31076 54068
rect 31128 53786 31156 54606
rect 30748 53780 30800 53786
rect 30748 53722 30800 53728
rect 31116 53780 31168 53786
rect 31116 53722 31168 53728
rect 31484 53712 31536 53718
rect 31484 53654 31536 53660
rect 31496 53242 31524 53654
rect 30472 53236 30524 53242
rect 30472 53178 30524 53184
rect 31484 53236 31536 53242
rect 31484 53178 31536 53184
rect 32048 52698 32076 57326
rect 32232 55146 32260 59200
rect 32588 57384 32640 57390
rect 32588 57326 32640 57332
rect 32312 56840 32364 56846
rect 32364 56800 32444 56828
rect 32312 56782 32364 56788
rect 32312 56704 32364 56710
rect 32312 56646 32364 56652
rect 32324 56370 32352 56646
rect 32312 56364 32364 56370
rect 32312 56306 32364 56312
rect 32416 55690 32444 56800
rect 32496 56160 32548 56166
rect 32496 56102 32548 56108
rect 32508 55894 32536 56102
rect 32496 55888 32548 55894
rect 32496 55830 32548 55836
rect 32600 55758 32628 57326
rect 32588 55752 32640 55758
rect 32588 55694 32640 55700
rect 32404 55684 32456 55690
rect 32404 55626 32456 55632
rect 32416 55282 32444 55626
rect 32404 55276 32456 55282
rect 32600 55264 32628 55694
rect 32692 55418 32720 59200
rect 32956 56840 33008 56846
rect 32956 56782 33008 56788
rect 32968 56710 32996 56782
rect 32956 56704 33008 56710
rect 32956 56646 33008 56652
rect 32968 56506 32996 56646
rect 32956 56500 33008 56506
rect 32956 56442 33008 56448
rect 32772 56364 32824 56370
rect 32772 56306 32824 56312
rect 32864 56364 32916 56370
rect 32864 56306 32916 56312
rect 32784 55826 32812 56306
rect 32772 55820 32824 55826
rect 32772 55762 32824 55768
rect 32876 55690 32904 56306
rect 33152 56250 33180 59200
rect 33416 57928 33468 57934
rect 33416 57870 33468 57876
rect 33428 56914 33456 57870
rect 33508 57452 33560 57458
rect 33508 57394 33560 57400
rect 33416 56908 33468 56914
rect 33416 56850 33468 56856
rect 33232 56840 33284 56846
rect 33232 56782 33284 56788
rect 33244 56438 33272 56782
rect 33520 56710 33548 57394
rect 33508 56704 33560 56710
rect 33508 56646 33560 56652
rect 33232 56432 33284 56438
rect 33232 56374 33284 56380
rect 33520 56370 33548 56646
rect 33508 56364 33560 56370
rect 33508 56306 33560 56312
rect 33152 56222 33364 56250
rect 33140 56160 33192 56166
rect 33140 56102 33192 56108
rect 33152 55758 33180 56102
rect 33140 55752 33192 55758
rect 33140 55694 33192 55700
rect 33232 55752 33284 55758
rect 33232 55694 33284 55700
rect 32864 55684 32916 55690
rect 32864 55626 32916 55632
rect 32680 55412 32732 55418
rect 32680 55354 32732 55360
rect 32680 55276 32732 55282
rect 32600 55236 32680 55264
rect 32404 55218 32456 55224
rect 32680 55218 32732 55224
rect 32220 55140 32272 55146
rect 32220 55082 32272 55088
rect 32128 54868 32180 54874
rect 32128 54810 32180 54816
rect 32140 53582 32168 54810
rect 32220 54528 32272 54534
rect 32220 54470 32272 54476
rect 32232 54126 32260 54470
rect 32220 54120 32272 54126
rect 32220 54062 32272 54068
rect 32232 53582 32260 54062
rect 32128 53576 32180 53582
rect 32128 53518 32180 53524
rect 32220 53576 32272 53582
rect 32220 53518 32272 53524
rect 32416 53242 32444 55218
rect 32588 54664 32640 54670
rect 32588 54606 32640 54612
rect 32496 54528 32548 54534
rect 32496 54470 32548 54476
rect 32508 54194 32536 54470
rect 32496 54188 32548 54194
rect 32496 54130 32548 54136
rect 32600 54126 32628 54606
rect 32692 54262 32720 55218
rect 33140 54664 33192 54670
rect 33140 54606 33192 54612
rect 32680 54256 32732 54262
rect 32680 54198 32732 54204
rect 32588 54120 32640 54126
rect 32588 54062 32640 54068
rect 33152 53786 33180 54606
rect 33244 54330 33272 55694
rect 33336 55282 33364 56222
rect 33612 56166 33640 59200
rect 33968 57792 34020 57798
rect 33968 57734 34020 57740
rect 33980 56982 34008 57734
rect 33968 56976 34020 56982
rect 33968 56918 34020 56924
rect 33968 56840 34020 56846
rect 33968 56782 34020 56788
rect 33600 56160 33652 56166
rect 33600 56102 33652 56108
rect 33980 55418 34008 56782
rect 34072 56234 34100 59200
rect 34532 57594 34560 59200
rect 34992 59106 35020 59200
rect 35084 59106 35112 59214
rect 34992 59078 35112 59106
rect 34520 57588 34572 57594
rect 34520 57530 34572 57536
rect 34244 57520 34296 57526
rect 34244 57462 34296 57468
rect 34152 57452 34204 57458
rect 34152 57394 34204 57400
rect 34164 56846 34192 57394
rect 34256 56846 34284 57462
rect 34336 57384 34388 57390
rect 34336 57326 34388 57332
rect 34152 56840 34204 56846
rect 34152 56782 34204 56788
rect 34244 56840 34296 56846
rect 34244 56782 34296 56788
rect 34164 56506 34192 56782
rect 34152 56500 34204 56506
rect 34152 56442 34204 56448
rect 34060 56228 34112 56234
rect 34060 56170 34112 56176
rect 34256 56001 34284 56782
rect 34348 56370 34376 57326
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 34888 56772 34940 56778
rect 34888 56714 34940 56720
rect 34336 56364 34388 56370
rect 34336 56306 34388 56312
rect 34242 55992 34298 56001
rect 34242 55927 34298 55936
rect 34256 55758 34284 55927
rect 34060 55752 34112 55758
rect 34060 55694 34112 55700
rect 34244 55752 34296 55758
rect 34244 55694 34296 55700
rect 34072 55593 34100 55694
rect 34058 55584 34114 55593
rect 34058 55519 34114 55528
rect 33784 55412 33836 55418
rect 33784 55354 33836 55360
rect 33968 55412 34020 55418
rect 33968 55354 34020 55360
rect 33324 55276 33376 55282
rect 33324 55218 33376 55224
rect 33796 55214 33824 55354
rect 33784 55208 33836 55214
rect 33784 55150 33836 55156
rect 33784 54868 33836 54874
rect 33784 54810 33836 54816
rect 33324 54596 33376 54602
rect 33324 54538 33376 54544
rect 33232 54324 33284 54330
rect 33232 54266 33284 54272
rect 33336 53990 33364 54538
rect 33324 53984 33376 53990
rect 33324 53926 33376 53932
rect 33140 53780 33192 53786
rect 33140 53722 33192 53728
rect 33336 53582 33364 53926
rect 33796 53786 33824 54810
rect 33968 54596 34020 54602
rect 33968 54538 34020 54544
rect 33784 53780 33836 53786
rect 33784 53722 33836 53728
rect 33324 53576 33376 53582
rect 33324 53518 33376 53524
rect 33796 53514 33824 53722
rect 33980 53650 34008 54538
rect 34072 54194 34100 55519
rect 34348 54602 34376 56306
rect 34704 56296 34756 56302
rect 34704 56238 34756 56244
rect 34428 56160 34480 56166
rect 34428 56102 34480 56108
rect 34440 55962 34468 56102
rect 34610 55992 34666 56001
rect 34428 55956 34480 55962
rect 34610 55927 34666 55936
rect 34428 55898 34480 55904
rect 34624 55758 34652 55927
rect 34716 55894 34744 56238
rect 34900 56234 34928 56714
rect 35360 56506 35388 59214
rect 35438 59200 35494 60000
rect 35898 59200 35954 60000
rect 36358 59200 36414 60000
rect 36818 59200 36874 60000
rect 37278 59200 37334 60000
rect 37738 59200 37794 60000
rect 38198 59200 38254 60000
rect 38658 59200 38714 60000
rect 39118 59200 39174 60000
rect 39578 59200 39634 60000
rect 40038 59200 40094 60000
rect 40144 59214 40356 59242
rect 35348 56500 35400 56506
rect 35348 56442 35400 56448
rect 34796 56228 34848 56234
rect 34796 56170 34848 56176
rect 34888 56228 34940 56234
rect 34888 56170 34940 56176
rect 34704 55888 34756 55894
rect 34704 55830 34756 55836
rect 34428 55752 34480 55758
rect 34428 55694 34480 55700
rect 34612 55752 34664 55758
rect 34612 55694 34664 55700
rect 34440 55604 34468 55694
rect 34440 55576 34652 55604
rect 34624 55418 34652 55576
rect 34612 55412 34664 55418
rect 34612 55354 34664 55360
rect 34520 55276 34572 55282
rect 34520 55218 34572 55224
rect 34336 54596 34388 54602
rect 34336 54538 34388 54544
rect 34336 54324 34388 54330
rect 34336 54266 34388 54272
rect 34060 54188 34112 54194
rect 34060 54130 34112 54136
rect 33968 53644 34020 53650
rect 33968 53586 34020 53592
rect 34072 53582 34100 54130
rect 34152 54120 34204 54126
rect 34152 54062 34204 54068
rect 34164 53582 34192 54062
rect 34348 53582 34376 54266
rect 34532 54262 34560 55218
rect 34704 55072 34756 55078
rect 34704 55014 34756 55020
rect 34520 54256 34572 54262
rect 34520 54198 34572 54204
rect 34716 54126 34744 55014
rect 34808 54874 34836 56170
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34888 55888 34940 55894
rect 34888 55830 34940 55836
rect 34900 55729 34928 55830
rect 35164 55820 35216 55826
rect 35164 55762 35216 55768
rect 34886 55720 34942 55729
rect 34886 55655 34942 55664
rect 35176 55418 35204 55762
rect 35348 55616 35400 55622
rect 35348 55558 35400 55564
rect 35164 55412 35216 55418
rect 35164 55354 35216 55360
rect 35360 55282 35388 55558
rect 35452 55350 35480 59200
rect 35912 57458 35940 59200
rect 35532 57452 35584 57458
rect 35532 57394 35584 57400
rect 35900 57452 35952 57458
rect 35900 57394 35952 57400
rect 35544 56914 35572 57394
rect 35716 57384 35768 57390
rect 35716 57326 35768 57332
rect 35532 56908 35584 56914
rect 35532 56850 35584 56856
rect 35728 56778 35756 57326
rect 35716 56772 35768 56778
rect 35716 56714 35768 56720
rect 35532 56432 35584 56438
rect 35532 56374 35584 56380
rect 35440 55344 35492 55350
rect 35440 55286 35492 55292
rect 35348 55276 35400 55282
rect 35348 55218 35400 55224
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34796 54868 34848 54874
rect 34796 54810 34848 54816
rect 35360 54194 35388 55218
rect 35544 55146 35572 56374
rect 35716 56364 35768 56370
rect 35716 56306 35768 56312
rect 35808 56364 35860 56370
rect 35808 56306 35860 56312
rect 35728 56234 35756 56306
rect 35716 56228 35768 56234
rect 35716 56170 35768 56176
rect 35624 56160 35676 56166
rect 35624 56102 35676 56108
rect 35636 55593 35664 56102
rect 35622 55584 35678 55593
rect 35622 55519 35678 55528
rect 35636 55282 35664 55519
rect 35624 55276 35676 55282
rect 35624 55218 35676 55224
rect 35532 55140 35584 55146
rect 35532 55082 35584 55088
rect 35544 54330 35572 55082
rect 35728 54806 35756 56170
rect 35820 54874 35848 56306
rect 35808 54868 35860 54874
rect 35808 54810 35860 54816
rect 35716 54800 35768 54806
rect 35716 54742 35768 54748
rect 35532 54324 35584 54330
rect 35532 54266 35584 54272
rect 35348 54188 35400 54194
rect 35348 54130 35400 54136
rect 34704 54120 34756 54126
rect 34704 54062 34756 54068
rect 34796 54120 34848 54126
rect 34796 54062 34848 54068
rect 34716 53650 34744 54062
rect 34808 53786 34836 54062
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 35544 53786 35572 54266
rect 35912 53786 35940 57394
rect 36268 57384 36320 57390
rect 36268 57326 36320 57332
rect 35992 56840 36044 56846
rect 35992 56782 36044 56788
rect 36004 56409 36032 56782
rect 36280 56438 36308 57326
rect 36268 56432 36320 56438
rect 35990 56400 36046 56409
rect 36268 56374 36320 56380
rect 35990 56335 36046 56344
rect 34796 53780 34848 53786
rect 34796 53722 34848 53728
rect 35532 53780 35584 53786
rect 35532 53722 35584 53728
rect 35900 53780 35952 53786
rect 35900 53722 35952 53728
rect 34704 53644 34756 53650
rect 34704 53586 34756 53592
rect 34060 53576 34112 53582
rect 34060 53518 34112 53524
rect 34152 53576 34204 53582
rect 34152 53518 34204 53524
rect 34336 53576 34388 53582
rect 34336 53518 34388 53524
rect 33784 53508 33836 53514
rect 33784 53450 33836 53456
rect 32404 53236 32456 53242
rect 32404 53178 32456 53184
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 32036 52692 32088 52698
rect 32036 52634 32088 52640
rect 36004 52086 36032 56335
rect 36372 55214 36400 59200
rect 36636 57384 36688 57390
rect 36636 57326 36688 57332
rect 36452 57044 36504 57050
rect 36452 56986 36504 56992
rect 36544 57044 36596 57050
rect 36544 56986 36596 56992
rect 36464 56438 36492 56986
rect 36556 56846 36584 56986
rect 36544 56840 36596 56846
rect 36544 56782 36596 56788
rect 36452 56432 36504 56438
rect 36452 56374 36504 56380
rect 36556 56370 36584 56782
rect 36544 56364 36596 56370
rect 36544 56306 36596 56312
rect 36648 55418 36676 57326
rect 36728 57316 36780 57322
rect 36728 57258 36780 57264
rect 36740 56846 36768 57258
rect 36832 56930 36860 59200
rect 37292 57458 37320 59200
rect 37280 57452 37332 57458
rect 37280 57394 37332 57400
rect 36832 56902 37044 56930
rect 36728 56840 36780 56846
rect 36728 56782 36780 56788
rect 36912 56840 36964 56846
rect 36912 56782 36964 56788
rect 36740 56438 36768 56782
rect 36728 56432 36780 56438
rect 36728 56374 36780 56380
rect 36924 56370 36952 56782
rect 36912 56364 36964 56370
rect 36912 56306 36964 56312
rect 36820 56160 36872 56166
rect 36820 56102 36872 56108
rect 36832 55826 36860 56102
rect 36924 55962 36952 56306
rect 36912 55956 36964 55962
rect 36912 55898 36964 55904
rect 36820 55820 36872 55826
rect 36820 55762 36872 55768
rect 36636 55412 36688 55418
rect 36636 55354 36688 55360
rect 37016 55282 37044 56902
rect 37004 55276 37056 55282
rect 37004 55218 37056 55224
rect 36360 55208 36412 55214
rect 36360 55150 36412 55156
rect 36452 54800 36504 54806
rect 36452 54742 36504 54748
rect 36464 54330 36492 54742
rect 37292 54330 37320 57394
rect 37752 56438 37780 59200
rect 37740 56432 37792 56438
rect 37740 56374 37792 56380
rect 37832 56160 37884 56166
rect 37832 56102 37884 56108
rect 37844 55962 37872 56102
rect 37832 55956 37884 55962
rect 37832 55898 37884 55904
rect 37372 55140 37424 55146
rect 37372 55082 37424 55088
rect 37384 54874 37412 55082
rect 37372 54868 37424 54874
rect 37372 54810 37424 54816
rect 37844 54806 37872 55898
rect 38212 55894 38240 59200
rect 38672 57458 38700 59200
rect 38660 57452 38712 57458
rect 38660 57394 38712 57400
rect 38936 57316 38988 57322
rect 38936 57258 38988 57264
rect 38752 57248 38804 57254
rect 38752 57190 38804 57196
rect 38474 56944 38530 56953
rect 38474 56879 38530 56888
rect 38660 56908 38712 56914
rect 38488 56846 38516 56879
rect 38660 56850 38712 56856
rect 38476 56840 38528 56846
rect 38476 56782 38528 56788
rect 38292 56296 38344 56302
rect 38292 56238 38344 56244
rect 38200 55888 38252 55894
rect 38200 55830 38252 55836
rect 38200 55752 38252 55758
rect 38200 55694 38252 55700
rect 38212 55282 38240 55694
rect 38304 55282 38332 56238
rect 38568 55752 38620 55758
rect 38568 55694 38620 55700
rect 38476 55616 38528 55622
rect 38476 55558 38528 55564
rect 38488 55418 38516 55558
rect 38476 55412 38528 55418
rect 38476 55354 38528 55360
rect 38488 55282 38516 55354
rect 38580 55282 38608 55694
rect 38200 55276 38252 55282
rect 38200 55218 38252 55224
rect 38292 55276 38344 55282
rect 38292 55218 38344 55224
rect 38476 55276 38528 55282
rect 38476 55218 38528 55224
rect 38568 55276 38620 55282
rect 38568 55218 38620 55224
rect 38212 54874 38240 55218
rect 38672 55214 38700 56850
rect 38764 56506 38792 57190
rect 38752 56500 38804 56506
rect 38752 56442 38804 56448
rect 38660 55208 38712 55214
rect 38660 55150 38712 55156
rect 38200 54868 38252 54874
rect 38200 54810 38252 54816
rect 37832 54800 37884 54806
rect 37832 54742 37884 54748
rect 38948 54330 38976 57258
rect 39132 56794 39160 59200
rect 39132 56766 39252 56794
rect 39120 56704 39172 56710
rect 39120 56646 39172 56652
rect 39132 56234 39160 56646
rect 39224 56438 39252 56766
rect 39212 56432 39264 56438
rect 39212 56374 39264 56380
rect 39212 56296 39264 56302
rect 39264 56256 39344 56284
rect 39212 56238 39264 56244
rect 39120 56228 39172 56234
rect 39120 56170 39172 56176
rect 39132 55962 39160 56170
rect 39120 55956 39172 55962
rect 39120 55898 39172 55904
rect 39316 55622 39344 56256
rect 39396 56228 39448 56234
rect 39396 56170 39448 56176
rect 39408 55690 39436 56170
rect 39396 55684 39448 55690
rect 39396 55626 39448 55632
rect 39304 55616 39356 55622
rect 39488 55616 39540 55622
rect 39304 55558 39356 55564
rect 39408 55564 39488 55570
rect 39408 55558 39540 55564
rect 39316 55350 39344 55558
rect 39408 55542 39528 55558
rect 39304 55344 39356 55350
rect 39304 55286 39356 55292
rect 39408 55282 39436 55542
rect 39396 55276 39448 55282
rect 39396 55218 39448 55224
rect 39488 55276 39540 55282
rect 39488 55218 39540 55224
rect 39408 54670 39436 55218
rect 39500 54738 39528 55218
rect 39488 54732 39540 54738
rect 39488 54674 39540 54680
rect 39396 54664 39448 54670
rect 39396 54606 39448 54612
rect 36452 54324 36504 54330
rect 36452 54266 36504 54272
rect 37280 54324 37332 54330
rect 37280 54266 37332 54272
rect 38936 54324 38988 54330
rect 38936 54266 38988 54272
rect 39592 54194 39620 59200
rect 40052 59106 40080 59200
rect 40144 59106 40172 59214
rect 40052 59078 40172 59106
rect 39856 57452 39908 57458
rect 39856 57394 39908 57400
rect 39580 54188 39632 54194
rect 39580 54130 39632 54136
rect 39868 53242 39896 57394
rect 40130 56944 40186 56953
rect 40130 56879 40132 56888
rect 40184 56879 40186 56888
rect 40132 56850 40184 56856
rect 40038 56808 40094 56817
rect 40038 56743 40094 56752
rect 40052 56710 40080 56743
rect 40040 56704 40092 56710
rect 40040 56646 40092 56652
rect 40144 56594 40172 56850
rect 40224 56840 40276 56846
rect 40224 56782 40276 56788
rect 40236 56710 40264 56782
rect 40224 56704 40276 56710
rect 40224 56646 40276 56652
rect 39960 56566 40172 56594
rect 39960 56522 39988 56566
rect 39960 56494 40080 56522
rect 40052 56438 40080 56494
rect 39948 56432 40000 56438
rect 39948 56374 40000 56380
rect 40040 56432 40092 56438
rect 40040 56374 40092 56380
rect 39960 55298 39988 56374
rect 40132 56364 40184 56370
rect 40132 56306 40184 56312
rect 40040 56296 40092 56302
rect 40040 56238 40092 56244
rect 40052 55418 40080 56238
rect 40144 55962 40172 56306
rect 40132 55956 40184 55962
rect 40132 55898 40184 55904
rect 40224 55684 40276 55690
rect 40224 55626 40276 55632
rect 40040 55412 40092 55418
rect 40040 55354 40092 55360
rect 39960 55270 40080 55298
rect 40236 55282 40264 55626
rect 39948 55208 40000 55214
rect 39948 55150 40000 55156
rect 39960 54126 39988 55150
rect 40052 54806 40080 55270
rect 40224 55276 40276 55282
rect 40224 55218 40276 55224
rect 40236 54874 40264 55218
rect 40224 54868 40276 54874
rect 40224 54810 40276 54816
rect 40040 54800 40092 54806
rect 40040 54742 40092 54748
rect 40328 54194 40356 59214
rect 40498 59200 40554 60000
rect 40958 59200 41014 60000
rect 41418 59200 41474 60000
rect 41878 59200 41934 60000
rect 42338 59200 42394 60000
rect 42798 59200 42854 60000
rect 43258 59200 43314 60000
rect 43718 59200 43774 60000
rect 44178 59200 44234 60000
rect 44638 59200 44694 60000
rect 45098 59200 45154 60000
rect 45558 59200 45614 60000
rect 46018 59200 46074 60000
rect 46478 59200 46534 60000
rect 46938 59200 46994 60000
rect 47398 59200 47454 60000
rect 47858 59200 47914 60000
rect 48318 59200 48374 60000
rect 48778 59200 48834 60000
rect 49238 59200 49294 60000
rect 49698 59200 49754 60000
rect 50158 59200 50214 60000
rect 50618 59200 50674 60000
rect 51078 59200 51134 60000
rect 51538 59200 51594 60000
rect 51998 59200 52054 60000
rect 52458 59200 52514 60000
rect 52918 59200 52974 60000
rect 53378 59200 53434 60000
rect 53838 59200 53894 60000
rect 54298 59200 54354 60000
rect 54758 59200 54814 60000
rect 55218 59200 55274 60000
rect 55678 59200 55734 60000
rect 56138 59200 56194 60000
rect 40512 57338 40540 59200
rect 40512 57310 40632 57338
rect 40500 57248 40552 57254
rect 40500 57190 40552 57196
rect 40512 56914 40540 57190
rect 40500 56908 40552 56914
rect 40500 56850 40552 56856
rect 40500 56364 40552 56370
rect 40500 56306 40552 56312
rect 40512 55962 40540 56306
rect 40604 56001 40632 57310
rect 40684 57316 40736 57322
rect 40684 57258 40736 57264
rect 40696 56914 40724 57258
rect 40684 56908 40736 56914
rect 40684 56850 40736 56856
rect 40972 56409 41000 59200
rect 41432 57866 41460 59200
rect 41420 57860 41472 57866
rect 41420 57802 41472 57808
rect 41052 57452 41104 57458
rect 41052 57394 41104 57400
rect 41064 57050 41092 57394
rect 41788 57384 41840 57390
rect 41788 57326 41840 57332
rect 41236 57316 41288 57322
rect 41236 57258 41288 57264
rect 41052 57044 41104 57050
rect 41052 56986 41104 56992
rect 41248 56710 41276 57258
rect 41800 56846 41828 57326
rect 41788 56840 41840 56846
rect 41788 56782 41840 56788
rect 41236 56704 41288 56710
rect 41236 56646 41288 56652
rect 40958 56400 41014 56409
rect 40958 56335 41014 56344
rect 40776 56296 40828 56302
rect 40774 56264 40776 56273
rect 40828 56264 40830 56273
rect 40774 56199 40830 56208
rect 40960 56160 41012 56166
rect 40960 56102 41012 56108
rect 40590 55992 40646 56001
rect 40500 55956 40552 55962
rect 40590 55927 40646 55936
rect 40500 55898 40552 55904
rect 40972 55894 41000 56102
rect 40960 55888 41012 55894
rect 40960 55830 41012 55836
rect 40408 55684 40460 55690
rect 40408 55626 40460 55632
rect 40420 55282 40448 55626
rect 40408 55276 40460 55282
rect 40408 55218 40460 55224
rect 41144 55072 41196 55078
rect 41144 55014 41196 55020
rect 40500 54868 40552 54874
rect 40500 54810 40552 54816
rect 40512 54330 40540 54810
rect 40500 54324 40552 54330
rect 40500 54266 40552 54272
rect 41156 54194 41184 55014
rect 41248 54874 41276 56646
rect 41892 56273 41920 59200
rect 42156 56840 42208 56846
rect 42156 56782 42208 56788
rect 42168 56506 42196 56782
rect 42156 56500 42208 56506
rect 42156 56442 42208 56448
rect 41972 56296 42024 56302
rect 41878 56264 41934 56273
rect 41972 56238 42024 56244
rect 41878 56199 41934 56208
rect 41420 56160 41472 56166
rect 41420 56102 41472 56108
rect 41788 56160 41840 56166
rect 41788 56102 41840 56108
rect 41432 55865 41460 56102
rect 41418 55856 41474 55865
rect 41418 55791 41474 55800
rect 41696 55276 41748 55282
rect 41696 55218 41748 55224
rect 41708 54874 41736 55218
rect 41236 54868 41288 54874
rect 41236 54810 41288 54816
rect 41696 54868 41748 54874
rect 41696 54810 41748 54816
rect 41236 54732 41288 54738
rect 41236 54674 41288 54680
rect 40316 54188 40368 54194
rect 40316 54130 40368 54136
rect 41144 54188 41196 54194
rect 41144 54130 41196 54136
rect 39948 54120 40000 54126
rect 39948 54062 40000 54068
rect 39960 53718 39988 54062
rect 40328 53786 40356 54130
rect 41248 54126 41276 54674
rect 41800 54330 41828 56102
rect 41880 55956 41932 55962
rect 41880 55898 41932 55904
rect 41892 55690 41920 55898
rect 41880 55684 41932 55690
rect 41880 55626 41932 55632
rect 41984 54330 42012 56238
rect 42352 55350 42380 59200
rect 42812 57458 42840 59200
rect 42892 57792 42944 57798
rect 42892 57734 42944 57740
rect 42800 57452 42852 57458
rect 42800 57394 42852 57400
rect 42904 57202 42932 57734
rect 42984 57384 43036 57390
rect 42984 57326 43036 57332
rect 42628 57174 42932 57202
rect 42628 56386 42656 57174
rect 42904 57050 42932 57174
rect 42708 57044 42760 57050
rect 42708 56986 42760 56992
rect 42892 57044 42944 57050
rect 42892 56986 42944 56992
rect 42720 56506 42748 56986
rect 42892 56704 42944 56710
rect 42892 56646 42944 56652
rect 42708 56500 42760 56506
rect 42708 56442 42760 56448
rect 42444 56358 42656 56386
rect 42720 56370 42748 56442
rect 42708 56364 42760 56370
rect 42444 56302 42472 56358
rect 42708 56306 42760 56312
rect 42432 56296 42484 56302
rect 42432 56238 42484 56244
rect 42524 56296 42576 56302
rect 42524 56238 42576 56244
rect 42536 55758 42564 56238
rect 42720 55962 42748 56306
rect 42708 55956 42760 55962
rect 42708 55898 42760 55904
rect 42904 55758 42932 56646
rect 42996 56148 43024 57326
rect 43272 57050 43300 59200
rect 43628 57384 43680 57390
rect 43628 57326 43680 57332
rect 43352 57248 43404 57254
rect 43352 57190 43404 57196
rect 43260 57044 43312 57050
rect 43260 56986 43312 56992
rect 43364 56914 43392 57190
rect 43352 56908 43404 56914
rect 43352 56850 43404 56856
rect 43076 56840 43128 56846
rect 43076 56782 43128 56788
rect 43088 56370 43116 56782
rect 43640 56370 43668 57326
rect 43732 56545 43760 59200
rect 44088 57452 44140 57458
rect 44088 57394 44140 57400
rect 43996 57384 44048 57390
rect 43996 57326 44048 57332
rect 44008 56846 44036 57326
rect 43996 56840 44048 56846
rect 43996 56782 44048 56788
rect 43718 56536 43774 56545
rect 44008 56506 44036 56782
rect 43718 56471 43774 56480
rect 43996 56500 44048 56506
rect 43996 56442 44048 56448
rect 43076 56364 43128 56370
rect 43076 56306 43128 56312
rect 43168 56364 43220 56370
rect 43168 56306 43220 56312
rect 43628 56364 43680 56370
rect 43628 56306 43680 56312
rect 43904 56364 43956 56370
rect 43904 56306 43956 56312
rect 43076 56160 43128 56166
rect 42996 56120 43076 56148
rect 43076 56102 43128 56108
rect 42524 55752 42576 55758
rect 42524 55694 42576 55700
rect 42892 55752 42944 55758
rect 42892 55694 42944 55700
rect 42904 55570 42932 55694
rect 42904 55542 43024 55570
rect 42798 55448 42854 55457
rect 42798 55383 42800 55392
rect 42852 55383 42854 55392
rect 42892 55412 42944 55418
rect 42800 55354 42852 55360
rect 42892 55354 42944 55360
rect 42340 55344 42392 55350
rect 42340 55286 42392 55292
rect 42904 55282 42932 55354
rect 42156 55276 42208 55282
rect 42156 55218 42208 55224
rect 42892 55276 42944 55282
rect 42892 55218 42944 55224
rect 42064 55072 42116 55078
rect 42064 55014 42116 55020
rect 42076 54670 42104 55014
rect 42064 54664 42116 54670
rect 42064 54606 42116 54612
rect 41788 54324 41840 54330
rect 41788 54266 41840 54272
rect 41972 54324 42024 54330
rect 41972 54266 42024 54272
rect 41236 54120 41288 54126
rect 41236 54062 41288 54068
rect 40316 53780 40368 53786
rect 40316 53722 40368 53728
rect 41984 53718 42012 54266
rect 42076 53786 42104 54606
rect 42168 54534 42196 55218
rect 42708 55072 42760 55078
rect 42708 55014 42760 55020
rect 42156 54528 42208 54534
rect 42156 54470 42208 54476
rect 42616 54528 42668 54534
rect 42616 54470 42668 54476
rect 42168 54262 42196 54470
rect 42156 54256 42208 54262
rect 42156 54198 42208 54204
rect 42628 54194 42656 54470
rect 42720 54330 42748 55014
rect 42800 54732 42852 54738
rect 42904 54720 42932 55218
rect 42852 54692 42932 54720
rect 42800 54674 42852 54680
rect 42708 54324 42760 54330
rect 42708 54266 42760 54272
rect 42616 54188 42668 54194
rect 42616 54130 42668 54136
rect 42064 53780 42116 53786
rect 42064 53722 42116 53728
rect 39948 53712 40000 53718
rect 39948 53654 40000 53660
rect 41972 53712 42024 53718
rect 41972 53654 42024 53660
rect 42628 53446 42656 54130
rect 42720 53786 42748 54266
rect 42996 54194 43024 55542
rect 43088 55146 43116 56102
rect 43180 55962 43208 56306
rect 43260 56296 43312 56302
rect 43260 56238 43312 56244
rect 43168 55956 43220 55962
rect 43168 55898 43220 55904
rect 43272 55282 43300 56238
rect 43442 55992 43498 56001
rect 43442 55927 43444 55936
rect 43496 55927 43498 55936
rect 43444 55898 43496 55904
rect 43640 55690 43668 56306
rect 43628 55684 43680 55690
rect 43628 55626 43680 55632
rect 43260 55276 43312 55282
rect 43260 55218 43312 55224
rect 43076 55140 43128 55146
rect 43076 55082 43128 55088
rect 43088 54738 43116 55082
rect 43272 54738 43300 55218
rect 43076 54732 43128 54738
rect 43076 54674 43128 54680
rect 43260 54732 43312 54738
rect 43260 54674 43312 54680
rect 42984 54188 43036 54194
rect 42984 54130 43036 54136
rect 42708 53780 42760 53786
rect 42708 53722 42760 53728
rect 42996 53514 43024 54130
rect 43088 54126 43116 54674
rect 43272 54194 43300 54674
rect 43916 54670 43944 56306
rect 43996 55752 44048 55758
rect 43996 55694 44048 55700
rect 44008 55418 44036 55694
rect 43996 55412 44048 55418
rect 43996 55354 44048 55360
rect 43904 54664 43956 54670
rect 43904 54606 43956 54612
rect 44008 54194 44036 55354
rect 44100 55350 44128 57394
rect 44088 55344 44140 55350
rect 44088 55286 44140 55292
rect 44192 55282 44220 59200
rect 44272 57452 44324 57458
rect 44456 57452 44508 57458
rect 44272 57394 44324 57400
rect 44376 57412 44456 57440
rect 44284 55457 44312 57394
rect 44376 56914 44404 57412
rect 44456 57394 44508 57400
rect 44364 56908 44416 56914
rect 44364 56850 44416 56856
rect 44364 56772 44416 56778
rect 44364 56714 44416 56720
rect 44376 55894 44404 56714
rect 44652 56234 44680 59200
rect 44916 57452 44968 57458
rect 44916 57394 44968 57400
rect 44928 56370 44956 57394
rect 45112 56982 45140 59200
rect 45572 57526 45600 59200
rect 45928 57860 45980 57866
rect 45928 57802 45980 57808
rect 45744 57588 45796 57594
rect 45744 57530 45796 57536
rect 45560 57520 45612 57526
rect 45560 57462 45612 57468
rect 45468 57248 45520 57254
rect 45468 57190 45520 57196
rect 45100 56976 45152 56982
rect 45100 56918 45152 56924
rect 45192 56840 45244 56846
rect 45192 56782 45244 56788
rect 45204 56409 45232 56782
rect 45376 56772 45428 56778
rect 45376 56714 45428 56720
rect 45388 56506 45416 56714
rect 45376 56500 45428 56506
rect 45376 56442 45428 56448
rect 45190 56400 45246 56409
rect 44916 56364 44968 56370
rect 45190 56335 45246 56344
rect 44916 56306 44968 56312
rect 44824 56296 44876 56302
rect 44824 56238 44876 56244
rect 44640 56228 44692 56234
rect 44640 56170 44692 56176
rect 44364 55888 44416 55894
rect 44364 55830 44416 55836
rect 44836 55758 44864 56238
rect 44824 55752 44876 55758
rect 44824 55694 44876 55700
rect 44928 55622 44956 56306
rect 45388 55758 45416 56442
rect 45480 56166 45508 57190
rect 45468 56160 45520 56166
rect 45468 56102 45520 56108
rect 45480 55894 45508 56102
rect 45468 55888 45520 55894
rect 45468 55830 45520 55836
rect 45376 55752 45428 55758
rect 45376 55694 45428 55700
rect 44916 55616 44968 55622
rect 44916 55558 44968 55564
rect 44270 55448 44326 55457
rect 45572 55418 45600 57462
rect 45756 57390 45784 57530
rect 45744 57384 45796 57390
rect 45744 57326 45796 57332
rect 45652 57316 45704 57322
rect 45652 57258 45704 57264
rect 45664 56438 45692 57258
rect 45652 56432 45704 56438
rect 45652 56374 45704 56380
rect 45664 55894 45692 56374
rect 45756 56370 45784 57326
rect 45940 56846 45968 57802
rect 46032 57050 46060 59200
rect 46388 57248 46440 57254
rect 46388 57190 46440 57196
rect 46020 57044 46072 57050
rect 46020 56986 46072 56992
rect 45928 56840 45980 56846
rect 45928 56782 45980 56788
rect 45744 56364 45796 56370
rect 45744 56306 45796 56312
rect 45744 56160 45796 56166
rect 45744 56102 45796 56108
rect 45652 55888 45704 55894
rect 45652 55830 45704 55836
rect 45756 55690 45784 56102
rect 45744 55684 45796 55690
rect 45744 55626 45796 55632
rect 44270 55383 44272 55392
rect 44324 55383 44326 55392
rect 45560 55412 45612 55418
rect 44272 55354 44324 55360
rect 45560 55354 45612 55360
rect 45940 55350 45968 56782
rect 46400 56273 46428 57190
rect 46492 56370 46520 59200
rect 46848 57792 46900 57798
rect 46848 57734 46900 57740
rect 46480 56364 46532 56370
rect 46480 56306 46532 56312
rect 46860 56302 46888 57734
rect 46952 57390 46980 59200
rect 47412 57458 47440 59200
rect 47400 57452 47452 57458
rect 47400 57394 47452 57400
rect 46940 57384 46992 57390
rect 46940 57326 46992 57332
rect 47032 57248 47084 57254
rect 47032 57190 47084 57196
rect 47044 56545 47072 57190
rect 47030 56536 47086 56545
rect 47030 56471 47086 56480
rect 47872 56370 47900 59200
rect 48332 56914 48360 59200
rect 48320 56908 48372 56914
rect 48320 56850 48372 56856
rect 48792 56370 48820 59200
rect 49252 56370 49280 59200
rect 49712 57458 49740 59200
rect 49700 57452 49752 57458
rect 49700 57394 49752 57400
rect 49712 56506 49740 57394
rect 50172 57050 50200 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 50632 57050 50660 59200
rect 51092 57458 51120 59200
rect 51080 57452 51132 57458
rect 51080 57394 51132 57400
rect 51448 57452 51500 57458
rect 51448 57394 51500 57400
rect 50160 57044 50212 57050
rect 50160 56986 50212 56992
rect 50620 57044 50672 57050
rect 50620 56986 50672 56992
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 51460 56506 51488 57394
rect 51552 57050 51580 59200
rect 51816 57248 51868 57254
rect 51816 57190 51868 57196
rect 51540 57044 51592 57050
rect 51540 56986 51592 56992
rect 49700 56500 49752 56506
rect 49700 56442 49752 56448
rect 51448 56500 51500 56506
rect 51448 56442 51500 56448
rect 47860 56364 47912 56370
rect 47860 56306 47912 56312
rect 48780 56364 48832 56370
rect 48780 56306 48832 56312
rect 49240 56364 49292 56370
rect 49240 56306 49292 56312
rect 46848 56296 46900 56302
rect 46386 56264 46442 56273
rect 46848 56238 46900 56244
rect 46386 56199 46442 56208
rect 46860 55962 46888 56238
rect 46848 55956 46900 55962
rect 46848 55898 46900 55904
rect 51828 55826 51856 57190
rect 52012 57050 52040 59200
rect 52472 57526 52500 59200
rect 52460 57520 52512 57526
rect 52460 57462 52512 57468
rect 52932 57050 52960 59200
rect 53012 57520 53064 57526
rect 53012 57462 53064 57468
rect 52000 57044 52052 57050
rect 52000 56986 52052 56992
rect 52920 57044 52972 57050
rect 52920 56986 52972 56992
rect 53024 56506 53052 57462
rect 53104 57248 53156 57254
rect 53104 57190 53156 57196
rect 53012 56500 53064 56506
rect 53012 56442 53064 56448
rect 51816 55820 51868 55826
rect 51816 55762 51868 55768
rect 46204 55616 46256 55622
rect 46204 55558 46256 55564
rect 45928 55344 45980 55350
rect 45928 55286 45980 55292
rect 46216 55282 46244 55558
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 44180 55276 44232 55282
rect 44180 55218 44232 55224
rect 46204 55276 46256 55282
rect 46204 55218 46256 55224
rect 53116 55214 53144 57190
rect 53392 57050 53420 59200
rect 53852 57458 53880 59200
rect 54116 57792 54168 57798
rect 54116 57734 54168 57740
rect 54128 57594 54156 57734
rect 54116 57588 54168 57594
rect 54116 57530 54168 57536
rect 54312 57458 54340 59200
rect 53840 57452 53892 57458
rect 53840 57394 53892 57400
rect 54300 57452 54352 57458
rect 54300 57394 54352 57400
rect 53852 57050 53880 57394
rect 53380 57044 53432 57050
rect 53380 56986 53432 56992
rect 53840 57044 53892 57050
rect 53840 56986 53892 56992
rect 54772 56506 54800 59200
rect 55232 57458 55260 59200
rect 55220 57452 55272 57458
rect 55220 57394 55272 57400
rect 55692 57390 55720 59200
rect 56152 57458 56180 59200
rect 55772 57452 55824 57458
rect 55772 57394 55824 57400
rect 56140 57452 56192 57458
rect 56140 57394 56192 57400
rect 55680 57384 55732 57390
rect 55680 57326 55732 57332
rect 55784 57050 55812 57394
rect 55772 57044 55824 57050
rect 55772 56986 55824 56992
rect 55496 56840 55548 56846
rect 55496 56782 55548 56788
rect 55508 56506 55536 56782
rect 54760 56500 54812 56506
rect 54760 56442 54812 56448
rect 55496 56500 55548 56506
rect 55496 56442 55548 56448
rect 53104 55208 53156 55214
rect 53104 55150 53156 55156
rect 44180 54732 44232 54738
rect 44180 54674 44232 54680
rect 44192 54330 44220 54674
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 44180 54324 44232 54330
rect 44180 54266 44232 54272
rect 43260 54188 43312 54194
rect 43260 54130 43312 54136
rect 43996 54188 44048 54194
rect 43996 54130 44048 54136
rect 43076 54120 43128 54126
rect 43076 54062 43128 54068
rect 42984 53508 43036 53514
rect 42984 53450 43036 53456
rect 42616 53440 42668 53446
rect 42616 53382 42668 53388
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 39856 53236 39908 53242
rect 39856 53178 39908 53184
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 35992 52080 36044 52086
rect 35992 52022 36044 52028
rect 34152 51944 34204 51950
rect 34152 51886 34204 51892
rect 35716 51944 35768 51950
rect 35716 51886 35768 51892
rect 34164 51610 34192 51886
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34152 51604 34204 51610
rect 34152 51546 34204 51552
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 27344 7200 27396 7206
rect 27344 7142 27396 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 27356 6866 27384 7142
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 25056 5778 25084 6054
rect 25240 5778 25268 6598
rect 26436 6322 26464 6734
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 26528 6322 26556 6598
rect 26424 6316 26476 6322
rect 26424 6258 26476 6264
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 25044 5772 25096 5778
rect 25044 5714 25096 5720
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25964 5772 26016 5778
rect 25964 5714 26016 5720
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 25320 5024 25372 5030
rect 25320 4966 25372 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7668 800 7696 2382
rect 8220 800 8248 2790
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 8588 800 8616 2518
rect 8956 800 8984 3470
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9324 800 9352 2382
rect 9692 800 9720 2790
rect 9968 800 9996 3470
rect 10232 2848 10284 2854
rect 10232 2790 10284 2796
rect 10244 800 10272 2790
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10520 800 10548 2518
rect 10796 800 10824 3470
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11072 800 11100 2790
rect 11348 800 11376 2790
rect 11624 800 11652 3470
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11900 800 11928 2314
rect 12176 800 12204 2382
rect 12452 800 12480 3470
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12728 800 12756 2790
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13004 800 13032 2382
rect 13280 800 13308 3470
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13556 800 13584 2790
rect 13820 2508 13872 2514
rect 13820 2450 13872 2456
rect 13832 800 13860 2450
rect 14108 800 14136 3470
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14384 800 14412 2926
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14660 800 14688 2790
rect 14936 800 14964 3470
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15212 800 15240 2518
rect 15488 800 15516 2790
rect 15764 800 15792 3470
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16040 800 16068 2382
rect 16316 800 16344 2926
rect 16592 800 16620 3470
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 800 16896 2790
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 17144 800 17172 2518
rect 17328 800 17356 3878
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 17604 800 17632 3470
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17868 2508 17920 2514
rect 17868 2450 17920 2456
rect 17880 800 17908 2450
rect 18156 800 18184 2790
rect 18432 800 18460 3470
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18708 800 18736 2790
rect 18972 2576 19024 2582
rect 18972 2518 19024 2524
rect 18984 800 19012 2518
rect 19260 800 19288 3470
rect 19444 1986 19472 3878
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20076 2916 20128 2922
rect 20076 2858 20128 2864
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19444 1958 19564 1986
rect 19536 800 19564 1958
rect 19996 1306 20024 2450
rect 19812 1278 20024 1306
rect 19812 800 19840 1278
rect 20088 800 20116 2858
rect 20364 800 20392 3878
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20640 800 20668 3470
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20916 800 20944 2926
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 21192 800 21220 2314
rect 21468 800 21496 4558
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 21744 800 21772 3538
rect 22020 800 22048 3878
rect 22296 800 22324 4558
rect 23492 4146 23520 4558
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 22836 3664 22888 3670
rect 22836 3606 22888 3612
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22572 800 22600 2858
rect 22848 800 22876 3606
rect 23124 800 23152 3946
rect 23492 3534 23520 4082
rect 23572 3596 23624 3602
rect 23572 3538 23624 3544
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23492 3074 23520 3470
rect 23308 3058 23520 3074
rect 23296 3052 23520 3058
rect 23348 3046 23520 3052
rect 23296 2994 23348 3000
rect 23308 2446 23336 2994
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23492 2650 23520 2926
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23584 2582 23612 3538
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23400 800 23428 2450
rect 23676 800 23704 4966
rect 23848 4752 23900 4758
rect 23848 4694 23900 4700
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23768 1494 23796 2994
rect 23860 2394 23888 4694
rect 24688 4146 24716 4966
rect 25332 4690 25360 4966
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 25320 4004 25372 4010
rect 25320 3946 25372 3952
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23952 3126 23980 3470
rect 24044 3194 24348 3210
rect 24032 3188 24348 3194
rect 24084 3182 24348 3188
rect 24032 3130 24084 3136
rect 23940 3120 23992 3126
rect 23940 3062 23992 3068
rect 24320 3058 24348 3182
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24044 2446 24072 2994
rect 24032 2440 24084 2446
rect 23860 2366 23980 2394
rect 24032 2382 24084 2388
rect 23756 1488 23808 1494
rect 23756 1430 23808 1436
rect 23952 800 23980 2366
rect 24216 1488 24268 1494
rect 24216 1430 24268 1436
rect 24228 800 24256 1430
rect 24504 800 24532 3674
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 24780 3058 24808 3402
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24596 2938 24624 2994
rect 24596 2910 24808 2938
rect 24584 2848 24636 2854
rect 24584 2790 24636 2796
rect 24596 2514 24624 2790
rect 24584 2508 24636 2514
rect 24584 2450 24636 2456
rect 24780 800 24808 2910
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24872 2650 24900 2790
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 25044 2304 25096 2310
rect 25044 2246 25096 2252
rect 25056 800 25084 2246
rect 25332 800 25360 3946
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 25780 3664 25832 3670
rect 25780 3606 25832 3612
rect 25596 2372 25648 2378
rect 25596 2314 25648 2320
rect 25608 800 25636 2314
rect 25700 1850 25728 3606
rect 25792 3194 25820 3606
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 25792 2446 25820 3130
rect 25884 2446 25912 3878
rect 25976 2938 26004 5714
rect 26436 4826 26464 6258
rect 27356 5302 27384 6598
rect 27540 6254 27568 7822
rect 27620 7744 27672 7750
rect 27620 7686 27672 7692
rect 27632 6866 27660 7686
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27528 6112 27580 6118
rect 27528 6054 27580 6060
rect 27540 5778 27568 6054
rect 28000 5846 28028 7142
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 27804 5772 27856 5778
rect 27804 5714 27856 5720
rect 27344 5296 27396 5302
rect 27344 5238 27396 5244
rect 27712 5160 27764 5166
rect 27712 5102 27764 5108
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 26424 4820 26476 4826
rect 26424 4762 26476 4768
rect 26884 4752 26936 4758
rect 26884 4694 26936 4700
rect 26148 4616 26200 4622
rect 26148 4558 26200 4564
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 26068 4010 26096 4422
rect 26160 4282 26188 4558
rect 26148 4276 26200 4282
rect 26148 4218 26200 4224
rect 26896 4146 26924 4694
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 26056 4004 26108 4010
rect 26056 3946 26108 3952
rect 25976 2910 26188 2938
rect 25780 2440 25832 2446
rect 25780 2382 25832 2388
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 25700 1822 25912 1850
rect 25884 800 25912 1822
rect 26160 800 26188 2910
rect 26436 800 26464 4014
rect 27356 3602 27384 4966
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 26700 3596 26752 3602
rect 26700 3538 26752 3544
rect 27344 3596 27396 3602
rect 27344 3538 27396 3544
rect 26712 800 26740 3538
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 26988 800 27016 2926
rect 27632 2802 27660 4626
rect 27264 2774 27660 2802
rect 27264 800 27292 2774
rect 27724 2666 27752 5102
rect 27540 2638 27752 2666
rect 27540 800 27568 2638
rect 27816 800 27844 5714
rect 27896 2916 27948 2922
rect 27896 2858 27948 2864
rect 27908 2378 27936 2858
rect 27896 2372 27948 2378
rect 27896 2314 27948 2320
rect 28092 800 28120 6802
rect 29012 6322 29040 8570
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 29380 6390 29408 7686
rect 29564 7478 29592 7686
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29840 6798 29868 8570
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 30104 8288 30156 8294
rect 30104 8230 30156 8236
rect 30116 7886 30144 8230
rect 30104 7880 30156 7886
rect 30104 7822 30156 7828
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 29840 6458 29868 6734
rect 30116 6730 30144 7822
rect 30104 6724 30156 6730
rect 30104 6666 30156 6672
rect 29828 6452 29880 6458
rect 29828 6394 29880 6400
rect 29368 6384 29420 6390
rect 29368 6326 29420 6332
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 29184 6248 29236 6254
rect 29184 6190 29236 6196
rect 29736 6248 29788 6254
rect 29736 6190 29788 6196
rect 29196 4826 29224 6190
rect 29460 6112 29512 6118
rect 29460 6054 29512 6060
rect 29472 5234 29500 6054
rect 29460 5228 29512 5234
rect 29460 5170 29512 5176
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 29184 4820 29236 4826
rect 29184 4762 29236 4768
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 28368 800 28396 4014
rect 29656 3738 29684 5102
rect 29644 3732 29696 3738
rect 29644 3674 29696 3680
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28540 2508 28592 2514
rect 28540 2450 28592 2456
rect 28552 1170 28580 2450
rect 28552 1142 28672 1170
rect 28644 800 28672 1142
rect 28920 800 28948 3538
rect 29000 3120 29052 3126
rect 29000 3062 29052 3068
rect 29012 2378 29040 3062
rect 29184 2984 29236 2990
rect 29184 2926 29236 2932
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29196 800 29224 2926
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29472 800 29500 2790
rect 29748 800 29776 6190
rect 29920 5704 29972 5710
rect 29920 5646 29972 5652
rect 29932 4690 29960 5646
rect 29920 4684 29972 4690
rect 29920 4626 29972 4632
rect 30116 3534 30144 6666
rect 30484 5778 30512 7822
rect 30668 5778 30696 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 31116 7744 31168 7750
rect 31116 7686 31168 7692
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 30472 5772 30524 5778
rect 30472 5714 30524 5720
rect 30656 5772 30708 5778
rect 30656 5714 30708 5720
rect 30380 5160 30432 5166
rect 30380 5102 30432 5108
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30012 3460 30064 3466
rect 30012 3402 30064 3408
rect 30024 800 30052 3402
rect 30104 2984 30156 2990
rect 30104 2926 30156 2932
rect 30116 2310 30144 2926
rect 30196 2848 30248 2854
rect 30392 2802 30420 5102
rect 30564 4684 30616 4690
rect 30564 4626 30616 4632
rect 30472 4548 30524 4554
rect 30472 4490 30524 4496
rect 30484 3738 30512 4490
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 30196 2790 30248 2796
rect 30208 2514 30236 2790
rect 30300 2774 30420 2802
rect 30196 2508 30248 2514
rect 30196 2450 30248 2456
rect 30104 2304 30156 2310
rect 30104 2246 30156 2252
rect 30300 800 30328 2774
rect 30576 800 30604 4626
rect 30760 3466 30788 7278
rect 31128 6866 31156 7686
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31668 6860 31720 6866
rect 31668 6802 31720 6808
rect 30932 6792 30984 6798
rect 30932 6734 30984 6740
rect 30944 6322 30972 6734
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 31392 5772 31444 5778
rect 31392 5714 31444 5720
rect 30840 4072 30892 4078
rect 30840 4014 30892 4020
rect 30748 3460 30800 3466
rect 30748 3402 30800 3408
rect 30852 800 30880 4014
rect 31116 2984 31168 2990
rect 31116 2926 31168 2932
rect 31128 800 31156 2926
rect 31404 800 31432 5714
rect 31680 800 31708 6802
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 32772 6452 32824 6458
rect 32772 6394 32824 6400
rect 32784 5710 32812 6394
rect 35360 6322 35388 6734
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 33876 6248 33928 6254
rect 33876 6190 33928 6196
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 32496 5160 32548 5166
rect 32496 5102 32548 5108
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 31956 800 31984 2926
rect 32232 800 32260 3538
rect 32508 800 32536 5102
rect 32680 4684 32732 4690
rect 32680 4626 32732 4632
rect 32692 2774 32720 4626
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 32692 2746 32812 2774
rect 32784 800 32812 2746
rect 33060 800 33088 4014
rect 33600 3596 33652 3602
rect 33600 3538 33652 3544
rect 33324 2508 33376 2514
rect 33324 2450 33376 2456
rect 33336 800 33364 2450
rect 33612 800 33640 3538
rect 33888 800 33916 6190
rect 35624 6180 35676 6186
rect 35624 6122 35676 6128
rect 34152 6112 34204 6118
rect 34152 6054 34204 6060
rect 33968 5568 34020 5574
rect 33968 5510 34020 5516
rect 33980 5302 34008 5510
rect 33968 5296 34020 5302
rect 33968 5238 34020 5244
rect 34164 5234 34192 6054
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35636 5914 35664 6122
rect 35624 5908 35676 5914
rect 35624 5850 35676 5856
rect 35348 5772 35400 5778
rect 35348 5714 35400 5720
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 34152 5228 34204 5234
rect 34152 5170 34204 5176
rect 34532 4690 34560 5646
rect 34704 5160 34756 5166
rect 34704 5102 34756 5108
rect 34520 4684 34572 4690
rect 34520 4626 34572 4632
rect 34612 4140 34664 4146
rect 34612 4082 34664 4088
rect 34152 3732 34204 3738
rect 34152 3674 34204 3680
rect 34164 800 34192 3674
rect 34624 3670 34652 4082
rect 34716 3738 34744 5102
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35360 4622 35388 5714
rect 35348 4616 35400 4622
rect 35348 4558 35400 4564
rect 35532 4616 35584 4622
rect 35532 4558 35584 4564
rect 35360 4146 35388 4558
rect 35348 4140 35400 4146
rect 35348 4082 35400 4088
rect 35544 4078 35572 4558
rect 35624 4140 35676 4146
rect 35624 4082 35676 4088
rect 35532 4072 35584 4078
rect 35532 4014 35584 4020
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34704 3732 34756 3738
rect 34704 3674 34756 3680
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34612 3460 34664 3466
rect 34612 3402 34664 3408
rect 34428 2984 34480 2990
rect 34428 2926 34480 2932
rect 34440 800 34468 2926
rect 34624 2650 34652 3402
rect 34796 3120 34848 3126
rect 34796 3062 34848 3068
rect 34704 3052 34756 3058
rect 34704 2994 34756 3000
rect 34612 2644 34664 2650
rect 34612 2586 34664 2592
rect 34716 2582 34744 2994
rect 34704 2576 34756 2582
rect 34704 2518 34756 2524
rect 34808 2378 34836 3062
rect 35346 2816 35402 2825
rect 34934 2748 35242 2757
rect 35346 2751 35402 2760
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34704 2372 34756 2378
rect 34704 2314 34756 2320
rect 34796 2372 34848 2378
rect 34796 2314 34848 2320
rect 34716 2106 34744 2314
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34704 2100 34756 2106
rect 34704 2042 34756 2048
rect 34704 1420 34756 1426
rect 34704 1362 34756 1368
rect 34716 800 34744 1362
rect 34992 800 35020 2246
rect 35360 1442 35388 2751
rect 35452 2514 35480 3878
rect 35532 3732 35584 3738
rect 35532 3674 35584 3680
rect 35440 2508 35492 2514
rect 35440 2450 35492 2456
rect 35268 1414 35388 1442
rect 35268 800 35296 1414
rect 35544 800 35572 3674
rect 35636 2446 35664 4082
rect 35624 2440 35676 2446
rect 35624 2382 35676 2388
rect 35728 1426 35756 51886
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 36268 5568 36320 5574
rect 36268 5510 36320 5516
rect 36280 5302 36308 5510
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 36268 5296 36320 5302
rect 36268 5238 36320 5244
rect 36452 5160 36504 5166
rect 36452 5102 36504 5108
rect 36464 4826 36492 5102
rect 36452 4820 36504 4826
rect 36452 4762 36504 4768
rect 36820 4616 36872 4622
rect 36820 4558 36872 4564
rect 35808 4004 35860 4010
rect 35808 3946 35860 3952
rect 35716 1420 35768 1426
rect 35716 1362 35768 1368
rect 35820 800 35848 3946
rect 36832 3602 36860 4558
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 37188 4004 37240 4010
rect 37188 3946 37240 3952
rect 36912 3664 36964 3670
rect 36912 3606 36964 3612
rect 36820 3596 36872 3602
rect 36820 3538 36872 3544
rect 36360 3392 36412 3398
rect 36924 3346 36952 3606
rect 36360 3334 36412 3340
rect 36084 2916 36136 2922
rect 36084 2858 36136 2864
rect 36096 800 36124 2858
rect 36372 800 36400 3334
rect 36648 3318 36952 3346
rect 36648 800 36676 3318
rect 36912 3188 36964 3194
rect 36912 3130 36964 3136
rect 36924 800 36952 3130
rect 37200 800 37228 3946
rect 37384 3534 37412 4082
rect 38292 3936 38344 3942
rect 38292 3878 38344 3884
rect 39396 3936 39448 3942
rect 39396 3878 39448 3884
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37384 3058 37412 3470
rect 37648 3460 37700 3466
rect 37648 3402 37700 3408
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 37476 2650 37504 2926
rect 37556 2848 37608 2854
rect 37556 2790 37608 2796
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 37568 2106 37596 2790
rect 37556 2100 37608 2106
rect 37556 2042 37608 2048
rect 37660 1442 37688 3402
rect 37740 2916 37792 2922
rect 37740 2858 37792 2864
rect 37476 1414 37688 1442
rect 37476 800 37504 1414
rect 37752 800 37780 2858
rect 38016 2508 38068 2514
rect 38016 2450 38068 2456
rect 38028 800 38056 2450
rect 38304 800 38332 3878
rect 39120 3664 39172 3670
rect 39120 3606 39172 3612
rect 38844 2984 38896 2990
rect 38844 2926 38896 2932
rect 38750 2816 38806 2825
rect 38750 2751 38806 2760
rect 38764 2650 38792 2751
rect 38752 2644 38804 2650
rect 38752 2586 38804 2592
rect 38568 2440 38620 2446
rect 38568 2382 38620 2388
rect 38580 800 38608 2382
rect 38856 800 38884 2926
rect 39132 800 39160 3606
rect 39408 800 39436 3878
rect 41052 3664 41104 3670
rect 41052 3606 41104 3612
rect 45192 3664 45244 3670
rect 45192 3606 45244 3612
rect 47124 3664 47176 3670
rect 47124 3606 47176 3612
rect 39948 3596 40000 3602
rect 39948 3538 40000 3544
rect 39672 2916 39724 2922
rect 39672 2858 39724 2864
rect 39684 800 39712 2858
rect 39960 800 39988 3538
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 40040 3392 40092 3398
rect 40040 3334 40092 3340
rect 40052 2650 40080 3334
rect 40040 2644 40092 2650
rect 40040 2586 40092 2592
rect 40224 2372 40276 2378
rect 40224 2314 40276 2320
rect 40236 800 40264 2314
rect 40512 800 40540 3470
rect 40776 2984 40828 2990
rect 40776 2926 40828 2932
rect 40788 800 40816 2926
rect 41064 800 41092 3606
rect 41880 3596 41932 3602
rect 41880 3538 41932 3544
rect 42984 3596 43036 3602
rect 42984 3538 43036 3544
rect 41604 2916 41656 2922
rect 41604 2858 41656 2864
rect 41420 2508 41472 2514
rect 41420 2450 41472 2456
rect 41432 1442 41460 2450
rect 41340 1414 41460 1442
rect 41340 800 41368 1414
rect 41616 800 41644 2858
rect 41892 800 41920 3538
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42156 2576 42208 2582
rect 42156 2518 42208 2524
rect 42168 800 42196 2518
rect 42444 800 42472 3470
rect 42708 3052 42760 3058
rect 42708 2994 42760 3000
rect 42720 800 42748 2994
rect 42996 800 43024 3538
rect 44364 3528 44416 3534
rect 44364 3470 44416 3476
rect 43260 2984 43312 2990
rect 43260 2926 43312 2932
rect 43272 800 43300 2926
rect 43812 2848 43864 2854
rect 43812 2790 43864 2796
rect 43536 2508 43588 2514
rect 43536 2450 43588 2456
rect 43548 800 43576 2450
rect 43824 800 43852 2790
rect 44088 2372 44140 2378
rect 44088 2314 44140 2320
rect 44100 800 44128 2314
rect 44376 800 44404 3470
rect 44916 2916 44968 2922
rect 44916 2858 44968 2864
rect 44640 2576 44692 2582
rect 44640 2518 44692 2524
rect 44652 800 44680 2518
rect 44928 800 44956 2858
rect 45204 800 45232 3606
rect 45744 3528 45796 3534
rect 45744 3470 45796 3476
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 45480 800 45508 2790
rect 45756 800 45784 3470
rect 46296 3460 46348 3466
rect 46296 3402 46348 3408
rect 46020 2440 46072 2446
rect 46020 2382 46072 2388
rect 46032 800 46060 2382
rect 46308 800 46336 3402
rect 46848 2848 46900 2854
rect 46848 2790 46900 2796
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 46584 800 46612 2450
rect 46860 800 46888 2790
rect 47136 800 47164 3606
rect 47952 3528 48004 3534
rect 47952 3470 48004 3476
rect 49056 3528 49108 3534
rect 49056 3470 49108 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 50988 3528 51040 3534
rect 50988 3470 51040 3476
rect 51540 3528 51592 3534
rect 51540 3470 51592 3476
rect 47676 2916 47728 2922
rect 47676 2858 47728 2864
rect 47400 2372 47452 2378
rect 47400 2314 47452 2320
rect 47412 800 47440 2314
rect 47688 800 47716 2858
rect 47964 800 47992 3470
rect 48780 2984 48832 2990
rect 48780 2926 48832 2932
rect 48228 2848 48280 2854
rect 48228 2790 48280 2796
rect 48240 800 48268 2790
rect 48504 2576 48556 2582
rect 48504 2518 48556 2524
rect 48516 800 48544 2518
rect 48792 800 48820 2926
rect 49068 800 49096 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 49608 2916 49660 2922
rect 49608 2858 49660 2864
rect 49332 2508 49384 2514
rect 49332 2450 49384 2456
rect 49344 800 49372 2450
rect 49620 800 49648 2858
rect 50160 2848 50212 2854
rect 50160 2790 50212 2796
rect 49884 2440 49936 2446
rect 49884 2382 49936 2388
rect 49896 800 49924 2382
rect 50172 800 50200 2790
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1850 50660 3470
rect 50712 2916 50764 2922
rect 50712 2858 50764 2864
rect 50448 1822 50660 1850
rect 50448 800 50476 1822
rect 50724 800 50752 2858
rect 51000 800 51028 3470
rect 51264 2372 51316 2378
rect 51264 2314 51316 2320
rect 51276 800 51304 2314
rect 51552 800 51580 3470
rect 52092 2848 52144 2854
rect 52092 2790 52144 2796
rect 51816 2576 51868 2582
rect 51816 2518 51868 2524
rect 51828 800 51856 2518
rect 52104 800 52132 2790
rect 52368 2508 52420 2514
rect 52368 2450 52420 2456
rect 52380 800 52408 2450
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
<< via2 >>
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 6090 57332 6092 57352
rect 6092 57332 6144 57352
rect 6144 57332 6146 57352
rect 6090 57296 6146 57332
rect 12346 57452 12402 57488
rect 12346 57432 12348 57452
rect 12348 57432 12400 57452
rect 12400 57432 12402 57452
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 23846 56752 23902 56808
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 25594 55800 25650 55856
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 27158 57296 27214 57352
rect 27526 57432 27582 57488
rect 27618 56208 27674 56264
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 29366 56364 29422 56400
rect 29366 56344 29368 56364
rect 29368 56344 29420 56364
rect 29420 56344 29422 56364
rect 30286 55684 30342 55720
rect 30286 55664 30288 55684
rect 30288 55664 30340 55684
rect 30340 55664 30342 55684
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 34242 55936 34298 55992
rect 34058 55528 34114 55584
rect 34610 55936 34666 55992
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34886 55664 34942 55720
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 35622 55528 35678 55584
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 35990 56344 36046 56400
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 38474 56888 38530 56944
rect 40130 56908 40186 56944
rect 40130 56888 40132 56908
rect 40132 56888 40184 56908
rect 40184 56888 40186 56908
rect 40038 56752 40094 56808
rect 40958 56344 41014 56400
rect 40774 56244 40776 56264
rect 40776 56244 40828 56264
rect 40828 56244 40830 56264
rect 40774 56208 40830 56244
rect 40590 55936 40646 55992
rect 41878 56208 41934 56264
rect 41418 55800 41474 55856
rect 43718 56480 43774 56536
rect 42798 55412 42854 55448
rect 42798 55392 42800 55412
rect 42800 55392 42852 55412
rect 42852 55392 42854 55412
rect 43442 55956 43498 55992
rect 43442 55936 43444 55956
rect 43444 55936 43496 55956
rect 43496 55936 43498 55956
rect 45190 56344 45246 56400
rect 44270 55412 44326 55448
rect 44270 55392 44272 55412
rect 44272 55392 44324 55412
rect 44324 55392 44326 55412
rect 47030 56480 47086 56536
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 46386 56208 46442 56264
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35346 2760 35402 2816
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 38750 2760 38806 2816
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 12341 57490 12407 57493
rect 27521 57490 27587 57493
rect 12341 57488 27587 57490
rect 12341 57432 12346 57488
rect 12402 57432 27526 57488
rect 27582 57432 27587 57488
rect 12341 57430 27587 57432
rect 12341 57427 12407 57430
rect 27521 57427 27587 57430
rect 6085 57354 6151 57357
rect 27153 57354 27219 57357
rect 6085 57352 27219 57354
rect 6085 57296 6090 57352
rect 6146 57296 27158 57352
rect 27214 57296 27219 57352
rect 6085 57294 27219 57296
rect 6085 57291 6151 57294
rect 27153 57291 27219 57294
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 38469 56946 38535 56949
rect 40125 56946 40191 56949
rect 38469 56944 40191 56946
rect 38469 56888 38474 56944
rect 38530 56888 40130 56944
rect 40186 56888 40191 56944
rect 38469 56886 40191 56888
rect 38469 56883 38535 56886
rect 40125 56883 40191 56886
rect 23841 56810 23907 56813
rect 40033 56810 40099 56813
rect 23841 56808 40099 56810
rect 23841 56752 23846 56808
rect 23902 56752 40038 56808
rect 40094 56752 40099 56808
rect 23841 56750 40099 56752
rect 23841 56747 23907 56750
rect 40033 56747 40099 56750
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 43713 56538 43779 56541
rect 47025 56538 47091 56541
rect 43713 56536 47091 56538
rect 43713 56480 43718 56536
rect 43774 56480 47030 56536
rect 47086 56480 47091 56536
rect 43713 56478 47091 56480
rect 43713 56475 43779 56478
rect 47025 56475 47091 56478
rect 29361 56402 29427 56405
rect 35985 56402 36051 56405
rect 29361 56400 36051 56402
rect 29361 56344 29366 56400
rect 29422 56344 35990 56400
rect 36046 56344 36051 56400
rect 29361 56342 36051 56344
rect 29361 56339 29427 56342
rect 35985 56339 36051 56342
rect 40953 56402 41019 56405
rect 45185 56402 45251 56405
rect 40953 56400 45251 56402
rect 40953 56344 40958 56400
rect 41014 56344 45190 56400
rect 45246 56344 45251 56400
rect 40953 56342 45251 56344
rect 40953 56339 41019 56342
rect 45185 56339 45251 56342
rect 27613 56266 27679 56269
rect 40769 56266 40835 56269
rect 27613 56264 40835 56266
rect 27613 56208 27618 56264
rect 27674 56208 40774 56264
rect 40830 56208 40835 56264
rect 27613 56206 40835 56208
rect 27613 56203 27679 56206
rect 40769 56203 40835 56206
rect 41873 56266 41939 56269
rect 46381 56266 46447 56269
rect 41873 56264 46447 56266
rect 41873 56208 41878 56264
rect 41934 56208 46386 56264
rect 46442 56208 46447 56264
rect 41873 56206 46447 56208
rect 41873 56203 41939 56206
rect 46381 56203 46447 56206
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 34237 55994 34303 55997
rect 34605 55994 34671 55997
rect 34237 55992 34671 55994
rect 34237 55936 34242 55992
rect 34298 55936 34610 55992
rect 34666 55936 34671 55992
rect 34237 55934 34671 55936
rect 34237 55931 34303 55934
rect 34605 55931 34671 55934
rect 40585 55994 40651 55997
rect 43437 55994 43503 55997
rect 40585 55992 43503 55994
rect 40585 55936 40590 55992
rect 40646 55936 43442 55992
rect 43498 55936 43503 55992
rect 40585 55934 43503 55936
rect 40585 55931 40651 55934
rect 43437 55931 43503 55934
rect 25589 55858 25655 55861
rect 41413 55858 41479 55861
rect 25589 55856 41479 55858
rect 25589 55800 25594 55856
rect 25650 55800 41418 55856
rect 41474 55800 41479 55856
rect 25589 55798 41479 55800
rect 25589 55795 25655 55798
rect 41413 55795 41479 55798
rect 30281 55722 30347 55725
rect 34881 55722 34947 55725
rect 30281 55720 34947 55722
rect 30281 55664 30286 55720
rect 30342 55664 34886 55720
rect 34942 55664 34947 55720
rect 30281 55662 34947 55664
rect 30281 55659 30347 55662
rect 34881 55659 34947 55662
rect 34053 55586 34119 55589
rect 35617 55586 35683 55589
rect 34053 55584 35683 55586
rect 34053 55528 34058 55584
rect 34114 55528 35622 55584
rect 35678 55528 35683 55584
rect 34053 55526 35683 55528
rect 34053 55523 34119 55526
rect 35617 55523 35683 55526
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 42793 55450 42859 55453
rect 44265 55450 44331 55453
rect 42793 55448 44331 55450
rect 42793 55392 42798 55448
rect 42854 55392 44270 55448
rect 44326 55392 44331 55448
rect 42793 55390 44331 55392
rect 42793 55387 42859 55390
rect 44265 55387 44331 55390
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 35341 2818 35407 2821
rect 38745 2818 38811 2821
rect 35341 2816 38811 2818
rect 35341 2760 35346 2816
rect 35402 2760 38750 2816
rect 38806 2760 38811 2816
rect 35341 2758 38811 2760
rect 35341 2755 35407 2758
rect 38745 2755 38811 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 27324 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1666464484
transform 1 0 23828 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1666464484
transform -1 0 33120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1666464484
transform 1 0 29532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1666464484
transform 1 0 26128 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1666464484
transform 1 0 24748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A_N
timestamp 1666464484
transform 1 0 37168 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__B
timestamp 1666464484
transform 1 0 36340 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B1
timestamp 1666464484
transform 1 0 29072 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A_N
timestamp 1666464484
transform 1 0 46736 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__B1
timestamp 1666464484
transform 1 0 42780 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__235__B1
timestamp 1666464484
transform -1 0 28060 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1666464484
transform 1 0 35512 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__B2
timestamp 1666464484
transform 1 0 37536 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__A2
timestamp 1666464484
transform -1 0 31648 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A
timestamp 1666464484
transform -1 0 39468 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__A2
timestamp 1666464484
transform -1 0 41492 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1666464484
transform -1 0 23460 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__A
timestamp 1666464484
transform 1 0 24380 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A2
timestamp 1666464484
transform 1 0 36616 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A2
timestamp 1666464484
transform -1 0 34040 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1666464484
transform 1 0 36064 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__A1
timestamp 1666464484
transform 1 0 41952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A
timestamp 1666464484
transform 1 0 24932 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A
timestamp 1666464484
transform 1 0 25024 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A1
timestamp 1666464484
transform -1 0 33488 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A
timestamp 1666464484
transform -1 0 32936 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__B1
timestamp 1666464484
transform 1 0 31188 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 1666464484
transform 1 0 31372 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1666464484
transform 1 0 40756 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A1
timestamp 1666464484
transform -1 0 40940 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A
timestamp 1666464484
transform 1 0 25760 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A
timestamp 1666464484
transform 1 0 26496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A
timestamp 1666464484
transform 1 0 26864 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__285__A2
timestamp 1666464484
transform 1 0 39468 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A2
timestamp 1666464484
transform -1 0 34592 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__A1
timestamp 1666464484
transform 1 0 30728 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__295__C1
timestamp 1666464484
transform 1 0 26128 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1666464484
transform -1 0 3496 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1666464484
transform -1 0 27876 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1666464484
transform -1 0 30636 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1666464484
transform -1 0 32292 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1666464484
transform -1 0 35972 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1666464484
transform -1 0 39560 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1666464484
transform -1 0 35972 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1666464484
transform -1 0 37628 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1666464484
transform -1 0 40020 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1666464484
transform -1 0 40296 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1666464484
transform -1 0 45816 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1666464484
transform -1 0 46368 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1666464484
transform -1 0 45080 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1666464484
transform -1 0 46368 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1666464484
transform -1 0 49864 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1666464484
transform -1 0 49864 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1666464484
transform -1 0 50324 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1666464484
transform -1 0 51612 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1666464484
transform -1 0 53084 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1666464484
transform -1 0 54464 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1666464484
transform -1 0 56304 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_A
timestamp 1666464484
transform 1 0 5888 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1666464484
transform 1 0 11040 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_0_11
timestamp 1666464484
transform 1 0 2116 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_0_19
timestamp 1666464484
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_0_29
timestamp 1666464484
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_0_37
timestamp 1666464484
transform 1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_0_45
timestamp 1666464484
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 5980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1666464484
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_0_57
timestamp 1666464484
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_75
timestamp 1666464484
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1666464484
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_85
timestamp 1666464484
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_96
timestamp 1666464484
transform 1 0 9936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_103
timestamp 1666464484
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1666464484
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_113
timestamp 1666464484
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_124
timestamp 1666464484
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_131
timestamp 1666464484
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1666464484
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_141
timestamp 1666464484
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_152
timestamp 1666464484
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_159
timestamp 1666464484
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1666464484
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_169
timestamp 1666464484
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_180
timestamp 1666464484
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_187
timestamp 1666464484
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1666464484
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_197
timestamp 1666464484
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_208
timestamp 1666464484
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_215
timestamp 1666464484
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1666464484
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_225
timestamp 1666464484
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_236
timestamp 1666464484
transform 1 0 22816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_243
timestamp 1666464484
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1666464484
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_0_253
timestamp 1666464484
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_264
timestamp 1666464484
transform 1 0 25392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_271
timestamp 1666464484
transform 1 0 26036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1666464484
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_281
timestamp 1666464484
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_306
timestamp 1666464484
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1666464484
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_332
timestamp 1666464484
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_337
timestamp 1666464484
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1666464484
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1666464484
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_370
timestamp 1666464484
transform 1 0 35144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_377
timestamp 1666464484
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_384
timestamp 1666464484
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1666464484
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_398
timestamp 1666464484
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_405
timestamp 1666464484
transform 1 0 38364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_412
timestamp 1666464484
transform 1 0 39008 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1666464484
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_426
timestamp 1666464484
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_433
timestamp 1666464484
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_440
timestamp 1666464484
transform 1 0 41584 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1666464484
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_454
timestamp 1666464484
transform 1 0 42872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_461
timestamp 1666464484
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_468
timestamp 1666464484
transform 1 0 44160 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1666464484
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_482
timestamp 1666464484
transform 1 0 45448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_489
timestamp 1666464484
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_496
timestamp 1666464484
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1666464484
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_510
timestamp 1666464484
transform 1 0 48024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_517
timestamp 1666464484
transform 1 0 48668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_524
timestamp 1666464484
transform 1 0 49312 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1666464484
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_538
timestamp 1666464484
transform 1 0 50600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_545
timestamp 1666464484
transform 1 0 51244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_552
timestamp 1666464484
transform 1 0 51888 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_561
timestamp 1666464484
transform 1 0 52716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_566
timestamp 1666464484
transform 1 0 53176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_573
timestamp 1666464484
transform 1 0 53820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_580
timestamp 1666464484
transform 1 0 54464 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_0_589
timestamp 1666464484
transform 1 0 55292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_0_597
timestamp 1666464484
transform 1 0 56028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_0_605
timestamp 1666464484
transform 1 0 56764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_613
timestamp 1666464484
transform 1 0 57500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1666464484
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_0_617
timestamp 1666464484
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_3
timestamp 1666464484
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_11
timestamp 1666464484
transform 1 0 2116 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_19
timestamp 1666464484
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_27
timestamp 1666464484
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_35
timestamp 1666464484
transform 1 0 4324 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_43
timestamp 1666464484
transform 1 0 5060 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_1_51
timestamp 1666464484
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1666464484
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_1_57
timestamp 1666464484
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_65
timestamp 1666464484
transform 1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_1_73
timestamp 1666464484
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp 1666464484
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_81
timestamp 1666464484
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1666464484
transform 1 0 8924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_89
timestamp 1666464484
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_96
timestamp 1666464484
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_103
timestamp 1666464484
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1666464484
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_1_113
timestamp 1666464484
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_1_124
timestamp 1666464484
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_131
timestamp 1666464484
transform 1 0 13156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_138
timestamp 1666464484
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_145
timestamp 1666464484
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_152
timestamp 1666464484
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_159
timestamp 1666464484
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1666464484
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_1_169
timestamp 1666464484
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_1_180
timestamp 1666464484
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_187
timestamp 1666464484
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_194
timestamp 1666464484
transform 1 0 18952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_201
timestamp 1666464484
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_208
timestamp 1666464484
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_215
timestamp 1666464484
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1666464484
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_225
timestamp 1666464484
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_232
timestamp 1666464484
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_239
timestamp 1666464484
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_246
timestamp 1666464484
transform 1 0 23736 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_253
timestamp 1666464484
transform 1 0 24380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1666464484
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_281
timestamp 1666464484
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_285
timestamp 1666464484
transform 1 0 27324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_287
timestamp 1666464484
transform 1 0 27508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_309
timestamp 1666464484
transform 1 0 29532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_334
timestamp 1666464484
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1666464484
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_360
timestamp 1666464484
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_385
timestamp 1666464484
transform 1 0 36524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_389
timestamp 1666464484
transform 1 0 36892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1666464484
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1666464484
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_398
timestamp 1666464484
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_405
timestamp 1666464484
transform 1 0 38364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_412
timestamp 1666464484
transform 1 0 39008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_419
timestamp 1666464484
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_426
timestamp 1666464484
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_433
timestamp 1666464484
transform 1 0 40940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_1_440
timestamp 1666464484
transform 1 0 41584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1666464484
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_454
timestamp 1666464484
transform 1 0 42872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_461
timestamp 1666464484
transform 1 0 43516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_468
timestamp 1666464484
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_475
timestamp 1666464484
transform 1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_482
timestamp 1666464484
transform 1 0 45448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_489
timestamp 1666464484
transform 1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_1_496
timestamp 1666464484
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_505
timestamp 1666464484
transform 1 0 47564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_510
timestamp 1666464484
transform 1 0 48024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_517
timestamp 1666464484
transform 1 0 48668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_524
timestamp 1666464484
transform 1 0 49312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_531
timestamp 1666464484
transform 1 0 49956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_538
timestamp 1666464484
transform 1 0 50600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_545
timestamp 1666464484
transform 1 0 51244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_1_552
timestamp 1666464484
transform 1 0 51888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_561
timestamp 1666464484
transform 1 0 52716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_1_566
timestamp 1666464484
transform 1 0 53176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_574
timestamp 1666464484
transform 1 0 53912 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_582
timestamp 1666464484
transform 1 0 54648 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_590
timestamp 1666464484
transform 1 0 55384 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_598
timestamp 1666464484
transform 1 0 56120 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_1_606
timestamp 1666464484
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1666464484
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_1_617
timestamp 1666464484
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_3
timestamp 1666464484
transform 1 0 1380 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_11
timestamp 1666464484
transform 1 0 2116 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_19
timestamp 1666464484
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1666464484
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_2_29
timestamp 1666464484
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_37
timestamp 1666464484
transform 1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_45
timestamp 1666464484
transform 1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_53
timestamp 1666464484
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_61
timestamp 1666464484
transform 1 0 6716 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_69
timestamp 1666464484
transform 1 0 7452 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_2_77
timestamp 1666464484
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 1666464484
transform 1 0 8556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1666464484
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1666464484
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_90
timestamp 1666464484
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_94
timestamp 1666464484
transform 1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_96
timestamp 1666464484
transform 1 0 9936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_100
timestamp 1666464484
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_104
timestamp 1666464484
transform 1 0 10672 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_109
timestamp 1666464484
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1666464484
transform 1 0 11500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_118
timestamp 1666464484
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_122
timestamp 1666464484
transform 1 0 12328 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_127
timestamp 1666464484
transform 1 0 12788 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_131
timestamp 1666464484
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_136
timestamp 1666464484
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1666464484
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_146
timestamp 1666464484
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_150
timestamp 1666464484
transform 1 0 14904 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_154
timestamp 1666464484
transform 1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_158
timestamp 1666464484
transform 1 0 15640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_163
timestamp 1666464484
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1666464484
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_172
timestamp 1666464484
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_176
timestamp 1666464484
transform 1 0 17296 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_180
timestamp 1666464484
transform 1 0 17664 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_187
timestamp 1666464484
transform 1 0 18308 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1666464484
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_2_197
timestamp 1666464484
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_2_208
timestamp 1666464484
transform 1 0 20240 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_215
timestamp 1666464484
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_222
timestamp 1666464484
transform 1 0 21528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_229
timestamp 1666464484
transform 1 0 22172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_236
timestamp 1666464484
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_243
timestamp 1666464484
transform 1 0 23460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1666464484
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_253
timestamp 1666464484
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_257
timestamp 1666464484
transform 1 0 24748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_259
timestamp 1666464484
transform 1 0 24932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_281
timestamp 1666464484
transform 1 0 26956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1666464484
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1666464484
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_314
timestamp 1666464484
transform 1 0 29992 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_2_321
timestamp 1666464484
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_329
timestamp 1666464484
transform 1 0 31372 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_352
timestamp 1666464484
transform 1 0 33488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_359
timestamp 1666464484
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1666464484
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1666464484
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_388
timestamp 1666464484
transform 1 0 36800 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_395
timestamp 1666464484
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_402
timestamp 1666464484
transform 1 0 38088 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_409
timestamp 1666464484
transform 1 0 38732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_416
timestamp 1666464484
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1666464484
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_426
timestamp 1666464484
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_433
timestamp 1666464484
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_440
timestamp 1666464484
transform 1 0 41584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_447
timestamp 1666464484
transform 1 0 42228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_454
timestamp 1666464484
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_461
timestamp 1666464484
transform 1 0 43516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_2_468
timestamp 1666464484
transform 1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1666464484
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_482
timestamp 1666464484
transform 1 0 45448 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_489
timestamp 1666464484
transform 1 0 46092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_496
timestamp 1666464484
transform 1 0 46736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_503
timestamp 1666464484
transform 1 0 47380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_510
timestamp 1666464484
transform 1 0 48024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_517
timestamp 1666464484
transform 1 0 48668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_521
timestamp 1666464484
transform 1 0 49036 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_525
timestamp 1666464484
transform 1 0 49404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_529
timestamp 1666464484
transform 1 0 49772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1666464484
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_533
timestamp 1666464484
transform 1 0 50140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_540
timestamp 1666464484
transform 1 0 50784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_547
timestamp 1666464484
transform 1 0 51428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_2_554
timestamp 1666464484
transform 1 0 52072 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_562
timestamp 1666464484
transform 1 0 52808 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_570
timestamp 1666464484
transform 1 0 53544 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_578
timestamp 1666464484
transform 1 0 54280 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_586
timestamp 1666464484
transform 1 0 55016 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_2_589
timestamp 1666464484
transform 1 0 55292 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_597
timestamp 1666464484
transform 1 0 56028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_605
timestamp 1666464484
transform 1 0 56764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_2_613
timestamp 1666464484
transform 1 0 57500 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_2_621
timestamp 1666464484
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_3_3
timestamp 1666464484
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_11
timestamp 1666464484
transform 1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_19
timestamp 1666464484
transform 1 0 2852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_27
timestamp 1666464484
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_35
timestamp 1666464484
transform 1 0 4324 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_43
timestamp 1666464484
transform 1 0 5060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_51
timestamp 1666464484
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1666464484
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_57
timestamp 1666464484
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_65
timestamp 1666464484
transform 1 0 7084 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_73
timestamp 1666464484
transform 1 0 7820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_81
timestamp 1666464484
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_89
timestamp 1666464484
transform 1 0 9292 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_97
timestamp 1666464484
transform 1 0 10028 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_105
timestamp 1666464484
transform 1 0 10764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1666464484
transform 1 0 11132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1666464484
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_113
timestamp 1666464484
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_121
timestamp 1666464484
transform 1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_129
timestamp 1666464484
transform 1 0 12972 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_137
timestamp 1666464484
transform 1 0 13708 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_145
timestamp 1666464484
transform 1 0 14444 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_153
timestamp 1666464484
transform 1 0 15180 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_161
timestamp 1666464484
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_165
timestamp 1666464484
transform 1 0 16284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1666464484
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_169
timestamp 1666464484
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_180
timestamp 1666464484
transform 1 0 17664 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_188
timestamp 1666464484
transform 1 0 18400 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_196
timestamp 1666464484
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_200
timestamp 1666464484
transform 1 0 19504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_204
timestamp 1666464484
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1666464484
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_213
timestamp 1666464484
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1666464484
transform 1 0 21068 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1666464484
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_225
timestamp 1666464484
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_232
timestamp 1666464484
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_239
timestamp 1666464484
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_246
timestamp 1666464484
transform 1 0 23736 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_253
timestamp 1666464484
transform 1 0 24380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_278
timestamp 1666464484
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_281
timestamp 1666464484
transform 1 0 26956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_285
timestamp 1666464484
transform 1 0 27324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_287
timestamp 1666464484
transform 1 0 27508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_309
timestamp 1666464484
transform 1 0 29532 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1666464484
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_337
timestamp 1666464484
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_341
timestamp 1666464484
transform 1 0 32476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_364
timestamp 1666464484
transform 1 0 34592 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_371
timestamp 1666464484
transform 1 0 35236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_378
timestamp 1666464484
transform 1 0 35880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_385
timestamp 1666464484
transform 1 0 36524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_389
timestamp 1666464484
transform 1 0 36892 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1666464484
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_393
timestamp 1666464484
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_398
timestamp 1666464484
transform 1 0 37720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_405
timestamp 1666464484
transform 1 0 38364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_412
timestamp 1666464484
transform 1 0 39008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_416
timestamp 1666464484
transform 1 0 39376 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_420
timestamp 1666464484
transform 1 0 39744 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_428
timestamp 1666464484
transform 1 0 40480 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_436
timestamp 1666464484
transform 1 0 41216 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_444
timestamp 1666464484
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_3_449
timestamp 1666464484
transform 1 0 42412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_457
timestamp 1666464484
transform 1 0 43148 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_465
timestamp 1666464484
transform 1 0 43884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_473
timestamp 1666464484
transform 1 0 44620 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_481
timestamp 1666464484
transform 1 0 45356 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_489
timestamp 1666464484
transform 1 0 46092 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_497
timestamp 1666464484
transform 1 0 46828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_501
timestamp 1666464484
transform 1 0 47196 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1666464484
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_505
timestamp 1666464484
transform 1 0 47564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_513
timestamp 1666464484
transform 1 0 48300 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_521
timestamp 1666464484
transform 1 0 49036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_529
timestamp 1666464484
transform 1 0 49772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_537
timestamp 1666464484
transform 1 0 50508 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_545
timestamp 1666464484
transform 1 0 51244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_553
timestamp 1666464484
transform 1 0 51980 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_557
timestamp 1666464484
transform 1 0 52348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1666464484
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_561
timestamp 1666464484
transform 1 0 52716 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_569
timestamp 1666464484
transform 1 0 53452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_577
timestamp 1666464484
transform 1 0 54188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_585
timestamp 1666464484
transform 1 0 54924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_593
timestamp 1666464484
transform 1 0 55660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_3_601
timestamp 1666464484
transform 1 0 56396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_609
timestamp 1666464484
transform 1 0 57132 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_613
timestamp 1666464484
transform 1 0 57500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1666464484
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_617
timestamp 1666464484
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_3
timestamp 1666464484
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_11
timestamp 1666464484
transform 1 0 2116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_19
timestamp 1666464484
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1666464484
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_29
timestamp 1666464484
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_37
timestamp 1666464484
transform 1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_45
timestamp 1666464484
transform 1 0 5244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_53
timestamp 1666464484
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_61
timestamp 1666464484
transform 1 0 6716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_69
timestamp 1666464484
transform 1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_77
timestamp 1666464484
transform 1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_81
timestamp 1666464484
transform 1 0 8556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1666464484
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_85
timestamp 1666464484
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_93
timestamp 1666464484
transform 1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_101
timestamp 1666464484
transform 1 0 10396 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_109
timestamp 1666464484
transform 1 0 11132 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_117
timestamp 1666464484
transform 1 0 11868 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_125
timestamp 1666464484
transform 1 0 12604 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_133
timestamp 1666464484
transform 1 0 13340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1666464484
transform 1 0 13708 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1666464484
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_141
timestamp 1666464484
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_149
timestamp 1666464484
transform 1 0 14812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_157
timestamp 1666464484
transform 1 0 15548 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_165
timestamp 1666464484
transform 1 0 16284 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_173
timestamp 1666464484
transform 1 0 17020 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_181
timestamp 1666464484
transform 1 0 17756 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_189
timestamp 1666464484
transform 1 0 18492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1666464484
transform 1 0 18860 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1666464484
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_197
timestamp 1666464484
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_205
timestamp 1666464484
transform 1 0 19964 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_213
timestamp 1666464484
transform 1 0 20700 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_221
timestamp 1666464484
transform 1 0 21436 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_225
timestamp 1666464484
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_229
timestamp 1666464484
transform 1 0 22172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_234
timestamp 1666464484
transform 1 0 22632 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_238
timestamp 1666464484
transform 1 0 23000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_243
timestamp 1666464484
transform 1 0 23460 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1666464484
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1666464484
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_255
timestamp 1666464484
transform 1 0 24564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_259
timestamp 1666464484
transform 1 0 24932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_266
timestamp 1666464484
transform 1 0 25576 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_273
timestamp 1666464484
transform 1 0 26220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_298
timestamp 1666464484
transform 1 0 28520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_302
timestamp 1666464484
transform 1 0 28888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_306
timestamp 1666464484
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_309
timestamp 1666464484
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_334
timestamp 1666464484
transform 1 0 31832 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_359
timestamp 1666464484
transform 1 0 34132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1666464484
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_365
timestamp 1666464484
transform 1 0 34684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_370
timestamp 1666464484
transform 1 0 35144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_377
timestamp 1666464484
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_384
timestamp 1666464484
transform 1 0 36432 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_4_391
timestamp 1666464484
transform 1 0 37076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_399
timestamp 1666464484
transform 1 0 37812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_407
timestamp 1666464484
transform 1 0 38548 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_415
timestamp 1666464484
transform 1 0 39284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1666464484
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_421
timestamp 1666464484
transform 1 0 39836 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_429
timestamp 1666464484
transform 1 0 40572 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_437
timestamp 1666464484
transform 1 0 41308 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_445
timestamp 1666464484
transform 1 0 42044 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_453
timestamp 1666464484
transform 1 0 42780 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_461
timestamp 1666464484
transform 1 0 43516 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_469
timestamp 1666464484
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_473
timestamp 1666464484
transform 1 0 44620 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1666464484
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_477
timestamp 1666464484
transform 1 0 44988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_485
timestamp 1666464484
transform 1 0 45724 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_493
timestamp 1666464484
transform 1 0 46460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_501
timestamp 1666464484
transform 1 0 47196 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_509
timestamp 1666464484
transform 1 0 47932 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_517
timestamp 1666464484
transform 1 0 48668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_525
timestamp 1666464484
transform 1 0 49404 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_529
timestamp 1666464484
transform 1 0 49772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1666464484
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_533
timestamp 1666464484
transform 1 0 50140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_541
timestamp 1666464484
transform 1 0 50876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_549
timestamp 1666464484
transform 1 0 51612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_557
timestamp 1666464484
transform 1 0 52348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_565
timestamp 1666464484
transform 1 0 53084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_573
timestamp 1666464484
transform 1 0 53820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_581
timestamp 1666464484
transform 1 0 54556 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_585
timestamp 1666464484
transform 1 0 54924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1666464484
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_589
timestamp 1666464484
transform 1 0 55292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_597
timestamp 1666464484
transform 1 0 56028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_605
timestamp 1666464484
transform 1 0 56764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_4_613
timestamp 1666464484
transform 1 0 57500 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_4_621
timestamp 1666464484
transform 1 0 58236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_5_3
timestamp 1666464484
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_11
timestamp 1666464484
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_19
timestamp 1666464484
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_27
timestamp 1666464484
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_35
timestamp 1666464484
transform 1 0 4324 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_43
timestamp 1666464484
transform 1 0 5060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_51
timestamp 1666464484
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1666464484
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_57
timestamp 1666464484
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_65
timestamp 1666464484
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_73
timestamp 1666464484
transform 1 0 7820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_81
timestamp 1666464484
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_89
timestamp 1666464484
transform 1 0 9292 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_97
timestamp 1666464484
transform 1 0 10028 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_105
timestamp 1666464484
transform 1 0 10764 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_109
timestamp 1666464484
transform 1 0 11132 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1666464484
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_113
timestamp 1666464484
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_121
timestamp 1666464484
transform 1 0 12236 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_129
timestamp 1666464484
transform 1 0 12972 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_137
timestamp 1666464484
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_145
timestamp 1666464484
transform 1 0 14444 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_153
timestamp 1666464484
transform 1 0 15180 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_161
timestamp 1666464484
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1666464484
transform 1 0 16284 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1666464484
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_169
timestamp 1666464484
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_177
timestamp 1666464484
transform 1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_185
timestamp 1666464484
transform 1 0 18124 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_193
timestamp 1666464484
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_201
timestamp 1666464484
transform 1 0 19596 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_209
timestamp 1666464484
transform 1 0 20332 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_217
timestamp 1666464484
transform 1 0 21068 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1666464484
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1666464484
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_225
timestamp 1666464484
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_233
timestamp 1666464484
transform 1 0 22540 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_241
timestamp 1666464484
transform 1 0 23276 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_245
timestamp 1666464484
transform 1 0 23644 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_249
timestamp 1666464484
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_253
timestamp 1666464484
transform 1 0 24380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_257
timestamp 1666464484
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_264
timestamp 1666464484
transform 1 0 25392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_271
timestamp 1666464484
transform 1 0 26036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1666464484
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1666464484
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_304
timestamp 1666464484
transform 1 0 29072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_329
timestamp 1666464484
transform 1 0 31372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_333
timestamp 1666464484
transform 1 0 31740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1666464484
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_337
timestamp 1666464484
transform 1 0 32108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_360
timestamp 1666464484
transform 1 0 34224 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_385
timestamp 1666464484
transform 1 0 36524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_389
timestamp 1666464484
transform 1 0 36892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1666464484
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_393
timestamp 1666464484
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_401
timestamp 1666464484
transform 1 0 37996 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_409
timestamp 1666464484
transform 1 0 38732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_417
timestamp 1666464484
transform 1 0 39468 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_425
timestamp 1666464484
transform 1 0 40204 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_433
timestamp 1666464484
transform 1 0 40940 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_441
timestamp 1666464484
transform 1 0 41676 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_445
timestamp 1666464484
transform 1 0 42044 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1666464484
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_449
timestamp 1666464484
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_457
timestamp 1666464484
transform 1 0 43148 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_465
timestamp 1666464484
transform 1 0 43884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_473
timestamp 1666464484
transform 1 0 44620 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_481
timestamp 1666464484
transform 1 0 45356 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_489
timestamp 1666464484
transform 1 0 46092 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_497
timestamp 1666464484
transform 1 0 46828 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_501
timestamp 1666464484
transform 1 0 47196 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1666464484
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_505
timestamp 1666464484
transform 1 0 47564 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_513
timestamp 1666464484
transform 1 0 48300 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_521
timestamp 1666464484
transform 1 0 49036 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_529
timestamp 1666464484
transform 1 0 49772 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_537
timestamp 1666464484
transform 1 0 50508 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_545
timestamp 1666464484
transform 1 0 51244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_553
timestamp 1666464484
transform 1 0 51980 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_557
timestamp 1666464484
transform 1 0 52348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1666464484
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_561
timestamp 1666464484
transform 1 0 52716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_569
timestamp 1666464484
transform 1 0 53452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_577
timestamp 1666464484
transform 1 0 54188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_585
timestamp 1666464484
transform 1 0 54924 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_593
timestamp 1666464484
transform 1 0 55660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_5_601
timestamp 1666464484
transform 1 0 56396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_5_609
timestamp 1666464484
transform 1 0 57132 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_613
timestamp 1666464484
transform 1 0 57500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1666464484
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_5_617
timestamp 1666464484
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_3
timestamp 1666464484
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_11
timestamp 1666464484
transform 1 0 2116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_19
timestamp 1666464484
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1666464484
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_29
timestamp 1666464484
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_37
timestamp 1666464484
transform 1 0 4508 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_45
timestamp 1666464484
transform 1 0 5244 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_53
timestamp 1666464484
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_61
timestamp 1666464484
transform 1 0 6716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_69
timestamp 1666464484
transform 1 0 7452 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_77
timestamp 1666464484
transform 1 0 8188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1666464484
transform 1 0 8556 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1666464484
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_85
timestamp 1666464484
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_93
timestamp 1666464484
transform 1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_101
timestamp 1666464484
transform 1 0 10396 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_109
timestamp 1666464484
transform 1 0 11132 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_117
timestamp 1666464484
transform 1 0 11868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_125
timestamp 1666464484
transform 1 0 12604 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_133
timestamp 1666464484
transform 1 0 13340 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_137
timestamp 1666464484
transform 1 0 13708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1666464484
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_141
timestamp 1666464484
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_149
timestamp 1666464484
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_157
timestamp 1666464484
transform 1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_165
timestamp 1666464484
transform 1 0 16284 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_173
timestamp 1666464484
transform 1 0 17020 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_181
timestamp 1666464484
transform 1 0 17756 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_189
timestamp 1666464484
transform 1 0 18492 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_193
timestamp 1666464484
transform 1 0 18860 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1666464484
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_197
timestamp 1666464484
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_205
timestamp 1666464484
transform 1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_213
timestamp 1666464484
transform 1 0 20700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_221
timestamp 1666464484
transform 1 0 21436 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_229
timestamp 1666464484
transform 1 0 22172 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_237
timestamp 1666464484
transform 1 0 22908 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_245
timestamp 1666464484
transform 1 0 23644 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_249
timestamp 1666464484
transform 1 0 24012 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1666464484
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_253
timestamp 1666464484
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_257
timestamp 1666464484
transform 1 0 24748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_259
timestamp 1666464484
transform 1 0 24932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_281
timestamp 1666464484
transform 1 0 26956 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1666464484
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1666464484
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_311
timestamp 1666464484
transform 1 0 29716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_315
timestamp 1666464484
transform 1 0 30084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_340
timestamp 1666464484
transform 1 0 32384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_350
timestamp 1666464484
transform 1 0 33304 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_357
timestamp 1666464484
transform 1 0 33948 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_361
timestamp 1666464484
transform 1 0 34316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1666464484
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1666464484
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_6_370
timestamp 1666464484
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_377
timestamp 1666464484
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_6_384
timestamp 1666464484
transform 1 0 36432 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_392
timestamp 1666464484
transform 1 0 37168 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_400
timestamp 1666464484
transform 1 0 37904 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_408
timestamp 1666464484
transform 1 0 38640 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_416
timestamp 1666464484
transform 1 0 39376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_6_421
timestamp 1666464484
transform 1 0 39836 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_429
timestamp 1666464484
transform 1 0 40572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_437
timestamp 1666464484
transform 1 0 41308 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_445
timestamp 1666464484
transform 1 0 42044 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_453
timestamp 1666464484
transform 1 0 42780 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_461
timestamp 1666464484
transform 1 0 43516 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_469
timestamp 1666464484
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_473
timestamp 1666464484
transform 1 0 44620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1666464484
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_477
timestamp 1666464484
transform 1 0 44988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_485
timestamp 1666464484
transform 1 0 45724 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_493
timestamp 1666464484
transform 1 0 46460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_501
timestamp 1666464484
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_509
timestamp 1666464484
transform 1 0 47932 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_517
timestamp 1666464484
transform 1 0 48668 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_525
timestamp 1666464484
transform 1 0 49404 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_529
timestamp 1666464484
transform 1 0 49772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1666464484
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_533
timestamp 1666464484
transform 1 0 50140 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_541
timestamp 1666464484
transform 1 0 50876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_549
timestamp 1666464484
transform 1 0 51612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_557
timestamp 1666464484
transform 1 0 52348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_565
timestamp 1666464484
transform 1 0 53084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_573
timestamp 1666464484
transform 1 0 53820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_581
timestamp 1666464484
transform 1 0 54556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_585
timestamp 1666464484
transform 1 0 54924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1666464484
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_6_589
timestamp 1666464484
transform 1 0 55292 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_597
timestamp 1666464484
transform 1 0 56028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_605
timestamp 1666464484
transform 1 0 56764 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_613
timestamp 1666464484
transform 1 0 57500 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_621
timestamp 1666464484
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_7_3
timestamp 1666464484
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_11
timestamp 1666464484
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_19
timestamp 1666464484
transform 1 0 2852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_27
timestamp 1666464484
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_35
timestamp 1666464484
transform 1 0 4324 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_43
timestamp 1666464484
transform 1 0 5060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_51
timestamp 1666464484
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1666464484
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_57
timestamp 1666464484
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_65
timestamp 1666464484
transform 1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_73
timestamp 1666464484
transform 1 0 7820 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_81
timestamp 1666464484
transform 1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_89
timestamp 1666464484
transform 1 0 9292 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_97
timestamp 1666464484
transform 1 0 10028 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_105
timestamp 1666464484
transform 1 0 10764 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_109
timestamp 1666464484
transform 1 0 11132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1666464484
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_113
timestamp 1666464484
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_121
timestamp 1666464484
transform 1 0 12236 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_129
timestamp 1666464484
transform 1 0 12972 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_137
timestamp 1666464484
transform 1 0 13708 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_145
timestamp 1666464484
transform 1 0 14444 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_153
timestamp 1666464484
transform 1 0 15180 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_161
timestamp 1666464484
transform 1 0 15916 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_165
timestamp 1666464484
transform 1 0 16284 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1666464484
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_169
timestamp 1666464484
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_177
timestamp 1666464484
transform 1 0 17388 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_185
timestamp 1666464484
transform 1 0 18124 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_193
timestamp 1666464484
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_201
timestamp 1666464484
transform 1 0 19596 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_209
timestamp 1666464484
transform 1 0 20332 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_217
timestamp 1666464484
transform 1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1666464484
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1666464484
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_225
timestamp 1666464484
transform 1 0 21804 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_233
timestamp 1666464484
transform 1 0 22540 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_241
timestamp 1666464484
transform 1 0 23276 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_249
timestamp 1666464484
transform 1 0 24012 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_257
timestamp 1666464484
transform 1 0 24748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_261
timestamp 1666464484
transform 1 0 25116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_263
timestamp 1666464484
transform 1 0 25300 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_267
timestamp 1666464484
transform 1 0 25668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1666464484
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_281
timestamp 1666464484
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_283
timestamp 1666464484
transform 1 0 27140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_290
timestamp 1666464484
transform 1 0 27784 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_301
timestamp 1666464484
transform 1 0 28796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_326
timestamp 1666464484
transform 1 0 31096 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_333
timestamp 1666464484
transform 1 0 31740 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1666464484
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_337
timestamp 1666464484
transform 1 0 32108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_7_342
timestamp 1666464484
transform 1 0 32568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_348
timestamp 1666464484
transform 1 0 33120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_7_373
timestamp 1666464484
transform 1 0 35420 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_381
timestamp 1666464484
transform 1 0 36156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_389
timestamp 1666464484
transform 1 0 36892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1666464484
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_393
timestamp 1666464484
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_401
timestamp 1666464484
transform 1 0 37996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_409
timestamp 1666464484
transform 1 0 38732 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_417
timestamp 1666464484
transform 1 0 39468 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_425
timestamp 1666464484
transform 1 0 40204 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_433
timestamp 1666464484
transform 1 0 40940 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_441
timestamp 1666464484
transform 1 0 41676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_445
timestamp 1666464484
transform 1 0 42044 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1666464484
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_449
timestamp 1666464484
transform 1 0 42412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_457
timestamp 1666464484
transform 1 0 43148 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_465
timestamp 1666464484
transform 1 0 43884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_473
timestamp 1666464484
transform 1 0 44620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_481
timestamp 1666464484
transform 1 0 45356 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_489
timestamp 1666464484
transform 1 0 46092 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_497
timestamp 1666464484
transform 1 0 46828 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_501
timestamp 1666464484
transform 1 0 47196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1666464484
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_505
timestamp 1666464484
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_513
timestamp 1666464484
transform 1 0 48300 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_521
timestamp 1666464484
transform 1 0 49036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_529
timestamp 1666464484
transform 1 0 49772 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_537
timestamp 1666464484
transform 1 0 50508 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_545
timestamp 1666464484
transform 1 0 51244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_553
timestamp 1666464484
transform 1 0 51980 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_557
timestamp 1666464484
transform 1 0 52348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1666464484
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_561
timestamp 1666464484
transform 1 0 52716 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_569
timestamp 1666464484
transform 1 0 53452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_577
timestamp 1666464484
transform 1 0 54188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_585
timestamp 1666464484
transform 1 0 54924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_593
timestamp 1666464484
transform 1 0 55660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_7_601
timestamp 1666464484
transform 1 0 56396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_609
timestamp 1666464484
transform 1 0 57132 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_613
timestamp 1666464484
transform 1 0 57500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1666464484
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_617
timestamp 1666464484
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_3
timestamp 1666464484
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_11
timestamp 1666464484
transform 1 0 2116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_19
timestamp 1666464484
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1666464484
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_29
timestamp 1666464484
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_37
timestamp 1666464484
transform 1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_45
timestamp 1666464484
transform 1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_53
timestamp 1666464484
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_61
timestamp 1666464484
transform 1 0 6716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_69
timestamp 1666464484
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_77
timestamp 1666464484
transform 1 0 8188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_81
timestamp 1666464484
transform 1 0 8556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1666464484
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_85
timestamp 1666464484
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_93
timestamp 1666464484
transform 1 0 9660 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_101
timestamp 1666464484
transform 1 0 10396 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_109
timestamp 1666464484
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_117
timestamp 1666464484
transform 1 0 11868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_125
timestamp 1666464484
transform 1 0 12604 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_133
timestamp 1666464484
transform 1 0 13340 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_137
timestamp 1666464484
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1666464484
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_141
timestamp 1666464484
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_149
timestamp 1666464484
transform 1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_157
timestamp 1666464484
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_165
timestamp 1666464484
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_173
timestamp 1666464484
transform 1 0 17020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_181
timestamp 1666464484
transform 1 0 17756 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_189
timestamp 1666464484
transform 1 0 18492 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_193
timestamp 1666464484
transform 1 0 18860 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1666464484
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_197
timestamp 1666464484
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_205
timestamp 1666464484
transform 1 0 19964 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_213
timestamp 1666464484
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_221
timestamp 1666464484
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_229
timestamp 1666464484
transform 1 0 22172 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_237
timestamp 1666464484
transform 1 0 22908 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_245
timestamp 1666464484
transform 1 0 23644 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_249
timestamp 1666464484
transform 1 0 24012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1666464484
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_8_253
timestamp 1666464484
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_259
timestamp 1666464484
transform 1 0 24932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_266
timestamp 1666464484
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_270
timestamp 1666464484
transform 1 0 25944 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_8_274
timestamp 1666464484
transform 1 0 26312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_281
timestamp 1666464484
transform 1 0 26956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1666464484
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1666464484
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_8_317
timestamp 1666464484
transform 1 0 30268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_321
timestamp 1666464484
transform 1 0 30636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_323
timestamp 1666464484
transform 1 0 30820 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_345
timestamp 1666464484
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_356
timestamp 1666464484
transform 1 0 33856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_365
timestamp 1666464484
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_373
timestamp 1666464484
transform 1 0 35420 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_381
timestamp 1666464484
transform 1 0 36156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_389
timestamp 1666464484
transform 1 0 36892 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_397
timestamp 1666464484
transform 1 0 37628 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_405
timestamp 1666464484
transform 1 0 38364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_413
timestamp 1666464484
transform 1 0 39100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_417
timestamp 1666464484
transform 1 0 39468 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1666464484
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_421
timestamp 1666464484
transform 1 0 39836 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_429
timestamp 1666464484
transform 1 0 40572 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_437
timestamp 1666464484
transform 1 0 41308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_445
timestamp 1666464484
transform 1 0 42044 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_453
timestamp 1666464484
transform 1 0 42780 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_461
timestamp 1666464484
transform 1 0 43516 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_469
timestamp 1666464484
transform 1 0 44252 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_473
timestamp 1666464484
transform 1 0 44620 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1666464484
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_477
timestamp 1666464484
transform 1 0 44988 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_485
timestamp 1666464484
transform 1 0 45724 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_493
timestamp 1666464484
transform 1 0 46460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_501
timestamp 1666464484
transform 1 0 47196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_509
timestamp 1666464484
transform 1 0 47932 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_517
timestamp 1666464484
transform 1 0 48668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_525
timestamp 1666464484
transform 1 0 49404 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_529
timestamp 1666464484
transform 1 0 49772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1666464484
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_533
timestamp 1666464484
transform 1 0 50140 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_541
timestamp 1666464484
transform 1 0 50876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_549
timestamp 1666464484
transform 1 0 51612 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_557
timestamp 1666464484
transform 1 0 52348 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_565
timestamp 1666464484
transform 1 0 53084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_573
timestamp 1666464484
transform 1 0 53820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_581
timestamp 1666464484
transform 1 0 54556 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_585
timestamp 1666464484
transform 1 0 54924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1666464484
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_8_589
timestamp 1666464484
transform 1 0 55292 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_597
timestamp 1666464484
transform 1 0 56028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_605
timestamp 1666464484
transform 1 0 56764 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_8_613
timestamp 1666464484
transform 1 0 57500 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_621
timestamp 1666464484
transform 1 0 58236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_9_3
timestamp 1666464484
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_11
timestamp 1666464484
transform 1 0 2116 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_19
timestamp 1666464484
transform 1 0 2852 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_27
timestamp 1666464484
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_35
timestamp 1666464484
transform 1 0 4324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_43
timestamp 1666464484
transform 1 0 5060 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_51
timestamp 1666464484
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1666464484
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_57
timestamp 1666464484
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_65
timestamp 1666464484
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_73
timestamp 1666464484
transform 1 0 7820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_81
timestamp 1666464484
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_89
timestamp 1666464484
transform 1 0 9292 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_97
timestamp 1666464484
transform 1 0 10028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_105
timestamp 1666464484
transform 1 0 10764 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1666464484
transform 1 0 11132 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1666464484
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_113
timestamp 1666464484
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_121
timestamp 1666464484
transform 1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_129
timestamp 1666464484
transform 1 0 12972 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_137
timestamp 1666464484
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_145
timestamp 1666464484
transform 1 0 14444 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_153
timestamp 1666464484
transform 1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_161
timestamp 1666464484
transform 1 0 15916 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_165
timestamp 1666464484
transform 1 0 16284 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1666464484
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_169
timestamp 1666464484
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_177
timestamp 1666464484
transform 1 0 17388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_185
timestamp 1666464484
transform 1 0 18124 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_193
timestamp 1666464484
transform 1 0 18860 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_201
timestamp 1666464484
transform 1 0 19596 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_209
timestamp 1666464484
transform 1 0 20332 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_217
timestamp 1666464484
transform 1 0 21068 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1666464484
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1666464484
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_225
timestamp 1666464484
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_233
timestamp 1666464484
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_241
timestamp 1666464484
transform 1 0 23276 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_249
timestamp 1666464484
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_257
timestamp 1666464484
transform 1 0 24748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_265
timestamp 1666464484
transform 1 0 25484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_273
timestamp 1666464484
transform 1 0 26220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_277
timestamp 1666464484
transform 1 0 26588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1666464484
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_281
timestamp 1666464484
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_288
timestamp 1666464484
transform 1 0 27600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_295
timestamp 1666464484
transform 1 0 28244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_299
timestamp 1666464484
transform 1 0 28612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_303
timestamp 1666464484
transform 1 0 28980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_9_328
timestamp 1666464484
transform 1 0 31280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_337
timestamp 1666464484
transform 1 0 32108 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_345
timestamp 1666464484
transform 1 0 32844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_353
timestamp 1666464484
transform 1 0 33580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_361
timestamp 1666464484
transform 1 0 34316 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_369
timestamp 1666464484
transform 1 0 35052 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_377
timestamp 1666464484
transform 1 0 35788 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_385
timestamp 1666464484
transform 1 0 36524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_389
timestamp 1666464484
transform 1 0 36892 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1666464484
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_393
timestamp 1666464484
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_401
timestamp 1666464484
transform 1 0 37996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_409
timestamp 1666464484
transform 1 0 38732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_417
timestamp 1666464484
transform 1 0 39468 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_425
timestamp 1666464484
transform 1 0 40204 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_433
timestamp 1666464484
transform 1 0 40940 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_441
timestamp 1666464484
transform 1 0 41676 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_445
timestamp 1666464484
transform 1 0 42044 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1666464484
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_449
timestamp 1666464484
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_457
timestamp 1666464484
transform 1 0 43148 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_465
timestamp 1666464484
transform 1 0 43884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_473
timestamp 1666464484
transform 1 0 44620 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_481
timestamp 1666464484
transform 1 0 45356 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_489
timestamp 1666464484
transform 1 0 46092 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_497
timestamp 1666464484
transform 1 0 46828 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_501
timestamp 1666464484
transform 1 0 47196 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1666464484
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_505
timestamp 1666464484
transform 1 0 47564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_513
timestamp 1666464484
transform 1 0 48300 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_521
timestamp 1666464484
transform 1 0 49036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_529
timestamp 1666464484
transform 1 0 49772 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_537
timestamp 1666464484
transform 1 0 50508 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_545
timestamp 1666464484
transform 1 0 51244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_553
timestamp 1666464484
transform 1 0 51980 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_557
timestamp 1666464484
transform 1 0 52348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1666464484
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_561
timestamp 1666464484
transform 1 0 52716 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_569
timestamp 1666464484
transform 1 0 53452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_577
timestamp 1666464484
transform 1 0 54188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_585
timestamp 1666464484
transform 1 0 54924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_593
timestamp 1666464484
transform 1 0 55660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_9_601
timestamp 1666464484
transform 1 0 56396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_609
timestamp 1666464484
transform 1 0 57132 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_613
timestamp 1666464484
transform 1 0 57500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1666464484
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_617
timestamp 1666464484
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_3
timestamp 1666464484
transform 1 0 1380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_11
timestamp 1666464484
transform 1 0 2116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_19
timestamp 1666464484
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1666464484
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_29
timestamp 1666464484
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_37
timestamp 1666464484
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_45
timestamp 1666464484
transform 1 0 5244 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_53
timestamp 1666464484
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_61
timestamp 1666464484
transform 1 0 6716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_69
timestamp 1666464484
transform 1 0 7452 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_77
timestamp 1666464484
transform 1 0 8188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_81
timestamp 1666464484
transform 1 0 8556 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1666464484
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_85
timestamp 1666464484
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_93
timestamp 1666464484
transform 1 0 9660 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_101
timestamp 1666464484
transform 1 0 10396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_109
timestamp 1666464484
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_117
timestamp 1666464484
transform 1 0 11868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_125
timestamp 1666464484
transform 1 0 12604 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_133
timestamp 1666464484
transform 1 0 13340 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_137
timestamp 1666464484
transform 1 0 13708 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1666464484
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_141
timestamp 1666464484
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_149
timestamp 1666464484
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_157
timestamp 1666464484
transform 1 0 15548 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_165
timestamp 1666464484
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_173
timestamp 1666464484
transform 1 0 17020 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_181
timestamp 1666464484
transform 1 0 17756 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_189
timestamp 1666464484
transform 1 0 18492 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_193
timestamp 1666464484
transform 1 0 18860 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1666464484
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_197
timestamp 1666464484
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_205
timestamp 1666464484
transform 1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_213
timestamp 1666464484
transform 1 0 20700 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_221
timestamp 1666464484
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_229
timestamp 1666464484
transform 1 0 22172 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_237
timestamp 1666464484
transform 1 0 22908 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_245
timestamp 1666464484
transform 1 0 23644 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_249
timestamp 1666464484
transform 1 0 24012 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1666464484
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_253
timestamp 1666464484
transform 1 0 24380 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_261
timestamp 1666464484
transform 1 0 25116 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_269
timestamp 1666464484
transform 1 0 25852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_277
timestamp 1666464484
transform 1 0 26588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_285
timestamp 1666464484
transform 1 0 27324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_289
timestamp 1666464484
transform 1 0 27692 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_293
timestamp 1666464484
transform 1 0 28060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_301
timestamp 1666464484
transform 1 0 28796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1666464484
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1666464484
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_10_314
timestamp 1666464484
transform 1 0 29992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_318
timestamp 1666464484
transform 1 0 30360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_10_322
timestamp 1666464484
transform 1 0 30728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_10_329
timestamp 1666464484
transform 1 0 31372 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_337
timestamp 1666464484
transform 1 0 32108 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_345
timestamp 1666464484
transform 1 0 32844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_353
timestamp 1666464484
transform 1 0 33580 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_361
timestamp 1666464484
transform 1 0 34316 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1666464484
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_365
timestamp 1666464484
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_373
timestamp 1666464484
transform 1 0 35420 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_381
timestamp 1666464484
transform 1 0 36156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_389
timestamp 1666464484
transform 1 0 36892 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_397
timestamp 1666464484
transform 1 0 37628 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_405
timestamp 1666464484
transform 1 0 38364 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_413
timestamp 1666464484
transform 1 0 39100 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_417
timestamp 1666464484
transform 1 0 39468 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1666464484
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_421
timestamp 1666464484
transform 1 0 39836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_429
timestamp 1666464484
transform 1 0 40572 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_437
timestamp 1666464484
transform 1 0 41308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_445
timestamp 1666464484
transform 1 0 42044 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_453
timestamp 1666464484
transform 1 0 42780 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_461
timestamp 1666464484
transform 1 0 43516 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_469
timestamp 1666464484
transform 1 0 44252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_473
timestamp 1666464484
transform 1 0 44620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1666464484
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_477
timestamp 1666464484
transform 1 0 44988 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_485
timestamp 1666464484
transform 1 0 45724 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_493
timestamp 1666464484
transform 1 0 46460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_501
timestamp 1666464484
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_509
timestamp 1666464484
transform 1 0 47932 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_517
timestamp 1666464484
transform 1 0 48668 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_525
timestamp 1666464484
transform 1 0 49404 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_529
timestamp 1666464484
transform 1 0 49772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1666464484
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_533
timestamp 1666464484
transform 1 0 50140 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_541
timestamp 1666464484
transform 1 0 50876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_549
timestamp 1666464484
transform 1 0 51612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_557
timestamp 1666464484
transform 1 0 52348 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_565
timestamp 1666464484
transform 1 0 53084 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_573
timestamp 1666464484
transform 1 0 53820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_581
timestamp 1666464484
transform 1 0 54556 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_585
timestamp 1666464484
transform 1 0 54924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1666464484
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_589
timestamp 1666464484
transform 1 0 55292 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_597
timestamp 1666464484
transform 1 0 56028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_605
timestamp 1666464484
transform 1 0 56764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_10_613
timestamp 1666464484
transform 1 0 57500 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_621
timestamp 1666464484
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_11_3
timestamp 1666464484
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_11
timestamp 1666464484
transform 1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_19
timestamp 1666464484
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_27
timestamp 1666464484
transform 1 0 3588 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_35
timestamp 1666464484
transform 1 0 4324 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_43
timestamp 1666464484
transform 1 0 5060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_51
timestamp 1666464484
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1666464484
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_57
timestamp 1666464484
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_65
timestamp 1666464484
transform 1 0 7084 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_73
timestamp 1666464484
transform 1 0 7820 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_81
timestamp 1666464484
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_89
timestamp 1666464484
transform 1 0 9292 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_97
timestamp 1666464484
transform 1 0 10028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_105
timestamp 1666464484
transform 1 0 10764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1666464484
transform 1 0 11132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1666464484
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_113
timestamp 1666464484
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_121
timestamp 1666464484
transform 1 0 12236 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_129
timestamp 1666464484
transform 1 0 12972 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_137
timestamp 1666464484
transform 1 0 13708 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_145
timestamp 1666464484
transform 1 0 14444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_153
timestamp 1666464484
transform 1 0 15180 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_161
timestamp 1666464484
transform 1 0 15916 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_165
timestamp 1666464484
transform 1 0 16284 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1666464484
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_169
timestamp 1666464484
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_177
timestamp 1666464484
transform 1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_185
timestamp 1666464484
transform 1 0 18124 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_193
timestamp 1666464484
transform 1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_201
timestamp 1666464484
transform 1 0 19596 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_209
timestamp 1666464484
transform 1 0 20332 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_217
timestamp 1666464484
transform 1 0 21068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1666464484
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1666464484
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_225
timestamp 1666464484
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_233
timestamp 1666464484
transform 1 0 22540 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_241
timestamp 1666464484
transform 1 0 23276 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_249
timestamp 1666464484
transform 1 0 24012 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_257
timestamp 1666464484
transform 1 0 24748 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_265
timestamp 1666464484
transform 1 0 25484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_273
timestamp 1666464484
transform 1 0 26220 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_277
timestamp 1666464484
transform 1 0 26588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1666464484
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_281
timestamp 1666464484
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_289
timestamp 1666464484
transform 1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_297
timestamp 1666464484
transform 1 0 28428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_305
timestamp 1666464484
transform 1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_11_311
timestamp 1666464484
transform 1 0 29716 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_322
timestamp 1666464484
transform 1 0 30728 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_330
timestamp 1666464484
transform 1 0 31464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_334
timestamp 1666464484
transform 1 0 31832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_11_337
timestamp 1666464484
transform 1 0 32108 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_345
timestamp 1666464484
transform 1 0 32844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_353
timestamp 1666464484
transform 1 0 33580 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_361
timestamp 1666464484
transform 1 0 34316 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_369
timestamp 1666464484
transform 1 0 35052 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_377
timestamp 1666464484
transform 1 0 35788 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_385
timestamp 1666464484
transform 1 0 36524 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_389
timestamp 1666464484
transform 1 0 36892 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1666464484
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_393
timestamp 1666464484
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_401
timestamp 1666464484
transform 1 0 37996 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_409
timestamp 1666464484
transform 1 0 38732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_417
timestamp 1666464484
transform 1 0 39468 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_425
timestamp 1666464484
transform 1 0 40204 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_433
timestamp 1666464484
transform 1 0 40940 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_441
timestamp 1666464484
transform 1 0 41676 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_445
timestamp 1666464484
transform 1 0 42044 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1666464484
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_449
timestamp 1666464484
transform 1 0 42412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_457
timestamp 1666464484
transform 1 0 43148 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_465
timestamp 1666464484
transform 1 0 43884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_473
timestamp 1666464484
transform 1 0 44620 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_481
timestamp 1666464484
transform 1 0 45356 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_489
timestamp 1666464484
transform 1 0 46092 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_497
timestamp 1666464484
transform 1 0 46828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_501
timestamp 1666464484
transform 1 0 47196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1666464484
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_505
timestamp 1666464484
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_513
timestamp 1666464484
transform 1 0 48300 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_521
timestamp 1666464484
transform 1 0 49036 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_529
timestamp 1666464484
transform 1 0 49772 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_537
timestamp 1666464484
transform 1 0 50508 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_545
timestamp 1666464484
transform 1 0 51244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_553
timestamp 1666464484
transform 1 0 51980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_557
timestamp 1666464484
transform 1 0 52348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1666464484
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_561
timestamp 1666464484
transform 1 0 52716 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_569
timestamp 1666464484
transform 1 0 53452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_577
timestamp 1666464484
transform 1 0 54188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_585
timestamp 1666464484
transform 1 0 54924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_593
timestamp 1666464484
transform 1 0 55660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_601
timestamp 1666464484
transform 1 0 56396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_609
timestamp 1666464484
transform 1 0 57132 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_613
timestamp 1666464484
transform 1 0 57500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1666464484
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_617
timestamp 1666464484
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_3
timestamp 1666464484
transform 1 0 1380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_11
timestamp 1666464484
transform 1 0 2116 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_19
timestamp 1666464484
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1666464484
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_29
timestamp 1666464484
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_37
timestamp 1666464484
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_45
timestamp 1666464484
transform 1 0 5244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_53
timestamp 1666464484
transform 1 0 5980 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_61
timestamp 1666464484
transform 1 0 6716 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_69
timestamp 1666464484
transform 1 0 7452 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_77
timestamp 1666464484
transform 1 0 8188 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_81
timestamp 1666464484
transform 1 0 8556 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1666464484
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_85
timestamp 1666464484
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_93
timestamp 1666464484
transform 1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_101
timestamp 1666464484
transform 1 0 10396 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_109
timestamp 1666464484
transform 1 0 11132 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_117
timestamp 1666464484
transform 1 0 11868 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_125
timestamp 1666464484
transform 1 0 12604 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_133
timestamp 1666464484
transform 1 0 13340 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_137
timestamp 1666464484
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1666464484
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_141
timestamp 1666464484
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_149
timestamp 1666464484
transform 1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_157
timestamp 1666464484
transform 1 0 15548 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_165
timestamp 1666464484
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_173
timestamp 1666464484
transform 1 0 17020 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_181
timestamp 1666464484
transform 1 0 17756 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_189
timestamp 1666464484
transform 1 0 18492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1666464484
transform 1 0 18860 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1666464484
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_197
timestamp 1666464484
transform 1 0 19228 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_205
timestamp 1666464484
transform 1 0 19964 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_213
timestamp 1666464484
transform 1 0 20700 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_221
timestamp 1666464484
transform 1 0 21436 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_229
timestamp 1666464484
transform 1 0 22172 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_237
timestamp 1666464484
transform 1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_245
timestamp 1666464484
transform 1 0 23644 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_249
timestamp 1666464484
transform 1 0 24012 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1666464484
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_253
timestamp 1666464484
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_261
timestamp 1666464484
transform 1 0 25116 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_269
timestamp 1666464484
transform 1 0 25852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_277
timestamp 1666464484
transform 1 0 26588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_285
timestamp 1666464484
transform 1 0 27324 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_293
timestamp 1666464484
transform 1 0 28060 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_301
timestamp 1666464484
transform 1 0 28796 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_305
timestamp 1666464484
transform 1 0 29164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1666464484
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_309
timestamp 1666464484
transform 1 0 29532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_317
timestamp 1666464484
transform 1 0 30268 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_325
timestamp 1666464484
transform 1 0 31004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_333
timestamp 1666464484
transform 1 0 31740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_341
timestamp 1666464484
transform 1 0 32476 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_349
timestamp 1666464484
transform 1 0 33212 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_357
timestamp 1666464484
transform 1 0 33948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_361
timestamp 1666464484
transform 1 0 34316 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1666464484
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_365
timestamp 1666464484
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_373
timestamp 1666464484
transform 1 0 35420 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_381
timestamp 1666464484
transform 1 0 36156 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_389
timestamp 1666464484
transform 1 0 36892 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_397
timestamp 1666464484
transform 1 0 37628 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_405
timestamp 1666464484
transform 1 0 38364 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_413
timestamp 1666464484
transform 1 0 39100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_417
timestamp 1666464484
transform 1 0 39468 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1666464484
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_421
timestamp 1666464484
transform 1 0 39836 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_429
timestamp 1666464484
transform 1 0 40572 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_437
timestamp 1666464484
transform 1 0 41308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_445
timestamp 1666464484
transform 1 0 42044 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_453
timestamp 1666464484
transform 1 0 42780 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_461
timestamp 1666464484
transform 1 0 43516 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_469
timestamp 1666464484
transform 1 0 44252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_473
timestamp 1666464484
transform 1 0 44620 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1666464484
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_477
timestamp 1666464484
transform 1 0 44988 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_485
timestamp 1666464484
transform 1 0 45724 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_493
timestamp 1666464484
transform 1 0 46460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_501
timestamp 1666464484
transform 1 0 47196 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_509
timestamp 1666464484
transform 1 0 47932 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_517
timestamp 1666464484
transform 1 0 48668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_525
timestamp 1666464484
transform 1 0 49404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_529
timestamp 1666464484
transform 1 0 49772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1666464484
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_533
timestamp 1666464484
transform 1 0 50140 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_541
timestamp 1666464484
transform 1 0 50876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_549
timestamp 1666464484
transform 1 0 51612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_557
timestamp 1666464484
transform 1 0 52348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_565
timestamp 1666464484
transform 1 0 53084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_573
timestamp 1666464484
transform 1 0 53820 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_581
timestamp 1666464484
transform 1 0 54556 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_585
timestamp 1666464484
transform 1 0 54924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1666464484
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_12_589
timestamp 1666464484
transform 1 0 55292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_597
timestamp 1666464484
transform 1 0 56028 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_605
timestamp 1666464484
transform 1 0 56764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_12_613
timestamp 1666464484
transform 1 0 57500 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_12_621
timestamp 1666464484
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_13_3
timestamp 1666464484
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_11
timestamp 1666464484
transform 1 0 2116 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_19
timestamp 1666464484
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_27
timestamp 1666464484
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_35
timestamp 1666464484
transform 1 0 4324 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_43
timestamp 1666464484
transform 1 0 5060 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_51
timestamp 1666464484
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1666464484
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_57
timestamp 1666464484
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_65
timestamp 1666464484
transform 1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_73
timestamp 1666464484
transform 1 0 7820 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_81
timestamp 1666464484
transform 1 0 8556 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_89
timestamp 1666464484
transform 1 0 9292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_97
timestamp 1666464484
transform 1 0 10028 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_105
timestamp 1666464484
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1666464484
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1666464484
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_113
timestamp 1666464484
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_121
timestamp 1666464484
transform 1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_129
timestamp 1666464484
transform 1 0 12972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_137
timestamp 1666464484
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_145
timestamp 1666464484
transform 1 0 14444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_153
timestamp 1666464484
transform 1 0 15180 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_161
timestamp 1666464484
transform 1 0 15916 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1666464484
transform 1 0 16284 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1666464484
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_169
timestamp 1666464484
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_177
timestamp 1666464484
transform 1 0 17388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_185
timestamp 1666464484
transform 1 0 18124 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_193
timestamp 1666464484
transform 1 0 18860 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_201
timestamp 1666464484
transform 1 0 19596 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_209
timestamp 1666464484
transform 1 0 20332 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_217
timestamp 1666464484
transform 1 0 21068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1666464484
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1666464484
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_225
timestamp 1666464484
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_233
timestamp 1666464484
transform 1 0 22540 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_241
timestamp 1666464484
transform 1 0 23276 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_249
timestamp 1666464484
transform 1 0 24012 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_257
timestamp 1666464484
transform 1 0 24748 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_265
timestamp 1666464484
transform 1 0 25484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_273
timestamp 1666464484
transform 1 0 26220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_277
timestamp 1666464484
transform 1 0 26588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1666464484
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_281
timestamp 1666464484
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_289
timestamp 1666464484
transform 1 0 27692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_297
timestamp 1666464484
transform 1 0 28428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_305
timestamp 1666464484
transform 1 0 29164 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_313
timestamp 1666464484
transform 1 0 29900 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_321
timestamp 1666464484
transform 1 0 30636 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_329
timestamp 1666464484
transform 1 0 31372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_333
timestamp 1666464484
transform 1 0 31740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1666464484
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_337
timestamp 1666464484
transform 1 0 32108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_345
timestamp 1666464484
transform 1 0 32844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_353
timestamp 1666464484
transform 1 0 33580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_361
timestamp 1666464484
transform 1 0 34316 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_369
timestamp 1666464484
transform 1 0 35052 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_377
timestamp 1666464484
transform 1 0 35788 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_385
timestamp 1666464484
transform 1 0 36524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_389
timestamp 1666464484
transform 1 0 36892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1666464484
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_393
timestamp 1666464484
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_401
timestamp 1666464484
transform 1 0 37996 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_409
timestamp 1666464484
transform 1 0 38732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_417
timestamp 1666464484
transform 1 0 39468 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_425
timestamp 1666464484
transform 1 0 40204 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_433
timestamp 1666464484
transform 1 0 40940 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_441
timestamp 1666464484
transform 1 0 41676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_445
timestamp 1666464484
transform 1 0 42044 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1666464484
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_449
timestamp 1666464484
transform 1 0 42412 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_457
timestamp 1666464484
transform 1 0 43148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_465
timestamp 1666464484
transform 1 0 43884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_473
timestamp 1666464484
transform 1 0 44620 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_481
timestamp 1666464484
transform 1 0 45356 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_489
timestamp 1666464484
transform 1 0 46092 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_497
timestamp 1666464484
transform 1 0 46828 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_501
timestamp 1666464484
transform 1 0 47196 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1666464484
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_505
timestamp 1666464484
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_513
timestamp 1666464484
transform 1 0 48300 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_521
timestamp 1666464484
transform 1 0 49036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_529
timestamp 1666464484
transform 1 0 49772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_537
timestamp 1666464484
transform 1 0 50508 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_545
timestamp 1666464484
transform 1 0 51244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_553
timestamp 1666464484
transform 1 0 51980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_557
timestamp 1666464484
transform 1 0 52348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1666464484
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_561
timestamp 1666464484
transform 1 0 52716 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_569
timestamp 1666464484
transform 1 0 53452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_577
timestamp 1666464484
transform 1 0 54188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_585
timestamp 1666464484
transform 1 0 54924 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_593
timestamp 1666464484
transform 1 0 55660 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_13_601
timestamp 1666464484
transform 1 0 56396 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_609
timestamp 1666464484
transform 1 0 57132 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_613
timestamp 1666464484
transform 1 0 57500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1666464484
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_13_617
timestamp 1666464484
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_3
timestamp 1666464484
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_11
timestamp 1666464484
transform 1 0 2116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_19
timestamp 1666464484
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1666464484
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_29
timestamp 1666464484
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_37
timestamp 1666464484
transform 1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_45
timestamp 1666464484
transform 1 0 5244 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_53
timestamp 1666464484
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_61
timestamp 1666464484
transform 1 0 6716 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_69
timestamp 1666464484
transform 1 0 7452 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_77
timestamp 1666464484
transform 1 0 8188 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_81
timestamp 1666464484
transform 1 0 8556 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1666464484
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_85
timestamp 1666464484
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_93
timestamp 1666464484
transform 1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_101
timestamp 1666464484
transform 1 0 10396 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_109
timestamp 1666464484
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_117
timestamp 1666464484
transform 1 0 11868 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_125
timestamp 1666464484
transform 1 0 12604 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_133
timestamp 1666464484
transform 1 0 13340 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_137
timestamp 1666464484
transform 1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1666464484
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_141
timestamp 1666464484
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_149
timestamp 1666464484
transform 1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_157
timestamp 1666464484
transform 1 0 15548 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_165
timestamp 1666464484
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_173
timestamp 1666464484
transform 1 0 17020 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_181
timestamp 1666464484
transform 1 0 17756 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_189
timestamp 1666464484
transform 1 0 18492 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1666464484
transform 1 0 18860 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1666464484
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_197
timestamp 1666464484
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_205
timestamp 1666464484
transform 1 0 19964 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_213
timestamp 1666464484
transform 1 0 20700 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_221
timestamp 1666464484
transform 1 0 21436 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_229
timestamp 1666464484
transform 1 0 22172 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_237
timestamp 1666464484
transform 1 0 22908 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_245
timestamp 1666464484
transform 1 0 23644 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_249
timestamp 1666464484
transform 1 0 24012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1666464484
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_253
timestamp 1666464484
transform 1 0 24380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_261
timestamp 1666464484
transform 1 0 25116 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_269
timestamp 1666464484
transform 1 0 25852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_277
timestamp 1666464484
transform 1 0 26588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_285
timestamp 1666464484
transform 1 0 27324 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_293
timestamp 1666464484
transform 1 0 28060 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_301
timestamp 1666464484
transform 1 0 28796 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_305
timestamp 1666464484
transform 1 0 29164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1666464484
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_309
timestamp 1666464484
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_317
timestamp 1666464484
transform 1 0 30268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_325
timestamp 1666464484
transform 1 0 31004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_333
timestamp 1666464484
transform 1 0 31740 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_341
timestamp 1666464484
transform 1 0 32476 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_349
timestamp 1666464484
transform 1 0 33212 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_357
timestamp 1666464484
transform 1 0 33948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_361
timestamp 1666464484
transform 1 0 34316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1666464484
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_365
timestamp 1666464484
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_373
timestamp 1666464484
transform 1 0 35420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_381
timestamp 1666464484
transform 1 0 36156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_389
timestamp 1666464484
transform 1 0 36892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_397
timestamp 1666464484
transform 1 0 37628 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_405
timestamp 1666464484
transform 1 0 38364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_413
timestamp 1666464484
transform 1 0 39100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_417
timestamp 1666464484
transform 1 0 39468 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1666464484
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_421
timestamp 1666464484
transform 1 0 39836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_429
timestamp 1666464484
transform 1 0 40572 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_437
timestamp 1666464484
transform 1 0 41308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_445
timestamp 1666464484
transform 1 0 42044 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_453
timestamp 1666464484
transform 1 0 42780 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_461
timestamp 1666464484
transform 1 0 43516 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_469
timestamp 1666464484
transform 1 0 44252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_473
timestamp 1666464484
transform 1 0 44620 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1666464484
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_477
timestamp 1666464484
transform 1 0 44988 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_485
timestamp 1666464484
transform 1 0 45724 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_493
timestamp 1666464484
transform 1 0 46460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_501
timestamp 1666464484
transform 1 0 47196 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_509
timestamp 1666464484
transform 1 0 47932 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_517
timestamp 1666464484
transform 1 0 48668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_525
timestamp 1666464484
transform 1 0 49404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_529
timestamp 1666464484
transform 1 0 49772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1666464484
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_533
timestamp 1666464484
transform 1 0 50140 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_541
timestamp 1666464484
transform 1 0 50876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_549
timestamp 1666464484
transform 1 0 51612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_557
timestamp 1666464484
transform 1 0 52348 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_565
timestamp 1666464484
transform 1 0 53084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_573
timestamp 1666464484
transform 1 0 53820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_581
timestamp 1666464484
transform 1 0 54556 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_585
timestamp 1666464484
transform 1 0 54924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1666464484
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_14_589
timestamp 1666464484
transform 1 0 55292 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_597
timestamp 1666464484
transform 1 0 56028 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_605
timestamp 1666464484
transform 1 0 56764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_613
timestamp 1666464484
transform 1 0 57500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_621
timestamp 1666464484
transform 1 0 58236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_15_3
timestamp 1666464484
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_11
timestamp 1666464484
transform 1 0 2116 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_19
timestamp 1666464484
transform 1 0 2852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_27
timestamp 1666464484
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_35
timestamp 1666464484
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_43
timestamp 1666464484
transform 1 0 5060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_51
timestamp 1666464484
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1666464484
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_57
timestamp 1666464484
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_65
timestamp 1666464484
transform 1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_73
timestamp 1666464484
transform 1 0 7820 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_81
timestamp 1666464484
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_89
timestamp 1666464484
transform 1 0 9292 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_97
timestamp 1666464484
transform 1 0 10028 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_105
timestamp 1666464484
transform 1 0 10764 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1666464484
transform 1 0 11132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1666464484
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_113
timestamp 1666464484
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_121
timestamp 1666464484
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_129
timestamp 1666464484
transform 1 0 12972 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_137
timestamp 1666464484
transform 1 0 13708 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_145
timestamp 1666464484
transform 1 0 14444 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_153
timestamp 1666464484
transform 1 0 15180 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_161
timestamp 1666464484
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_165
timestamp 1666464484
transform 1 0 16284 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1666464484
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_169
timestamp 1666464484
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_177
timestamp 1666464484
transform 1 0 17388 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_185
timestamp 1666464484
transform 1 0 18124 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_193
timestamp 1666464484
transform 1 0 18860 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_201
timestamp 1666464484
transform 1 0 19596 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_209
timestamp 1666464484
transform 1 0 20332 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_217
timestamp 1666464484
transform 1 0 21068 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1666464484
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1666464484
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_225
timestamp 1666464484
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_233
timestamp 1666464484
transform 1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_241
timestamp 1666464484
transform 1 0 23276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_249
timestamp 1666464484
transform 1 0 24012 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_257
timestamp 1666464484
transform 1 0 24748 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_265
timestamp 1666464484
transform 1 0 25484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_273
timestamp 1666464484
transform 1 0 26220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_277
timestamp 1666464484
transform 1 0 26588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1666464484
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_281
timestamp 1666464484
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_289
timestamp 1666464484
transform 1 0 27692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_297
timestamp 1666464484
transform 1 0 28428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_305
timestamp 1666464484
transform 1 0 29164 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_313
timestamp 1666464484
transform 1 0 29900 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_321
timestamp 1666464484
transform 1 0 30636 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_329
timestamp 1666464484
transform 1 0 31372 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_333
timestamp 1666464484
transform 1 0 31740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1666464484
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_337
timestamp 1666464484
transform 1 0 32108 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_345
timestamp 1666464484
transform 1 0 32844 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_353
timestamp 1666464484
transform 1 0 33580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_361
timestamp 1666464484
transform 1 0 34316 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_369
timestamp 1666464484
transform 1 0 35052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_377
timestamp 1666464484
transform 1 0 35788 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_385
timestamp 1666464484
transform 1 0 36524 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_389
timestamp 1666464484
transform 1 0 36892 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1666464484
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_393
timestamp 1666464484
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_401
timestamp 1666464484
transform 1 0 37996 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_409
timestamp 1666464484
transform 1 0 38732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_417
timestamp 1666464484
transform 1 0 39468 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_425
timestamp 1666464484
transform 1 0 40204 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_433
timestamp 1666464484
transform 1 0 40940 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_441
timestamp 1666464484
transform 1 0 41676 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_445
timestamp 1666464484
transform 1 0 42044 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1666464484
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_449
timestamp 1666464484
transform 1 0 42412 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_457
timestamp 1666464484
transform 1 0 43148 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_465
timestamp 1666464484
transform 1 0 43884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_473
timestamp 1666464484
transform 1 0 44620 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_481
timestamp 1666464484
transform 1 0 45356 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_489
timestamp 1666464484
transform 1 0 46092 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_497
timestamp 1666464484
transform 1 0 46828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_501
timestamp 1666464484
transform 1 0 47196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1666464484
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_505
timestamp 1666464484
transform 1 0 47564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_513
timestamp 1666464484
transform 1 0 48300 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_521
timestamp 1666464484
transform 1 0 49036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_529
timestamp 1666464484
transform 1 0 49772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_537
timestamp 1666464484
transform 1 0 50508 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_545
timestamp 1666464484
transform 1 0 51244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_553
timestamp 1666464484
transform 1 0 51980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_557
timestamp 1666464484
transform 1 0 52348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1666464484
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_561
timestamp 1666464484
transform 1 0 52716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_569
timestamp 1666464484
transform 1 0 53452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_577
timestamp 1666464484
transform 1 0 54188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_585
timestamp 1666464484
transform 1 0 54924 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_593
timestamp 1666464484
transform 1 0 55660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_15_601
timestamp 1666464484
transform 1 0 56396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_609
timestamp 1666464484
transform 1 0 57132 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_613
timestamp 1666464484
transform 1 0 57500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1666464484
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_617
timestamp 1666464484
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_3
timestamp 1666464484
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_11
timestamp 1666464484
transform 1 0 2116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_19
timestamp 1666464484
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1666464484
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_29
timestamp 1666464484
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_37
timestamp 1666464484
transform 1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_45
timestamp 1666464484
transform 1 0 5244 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_53
timestamp 1666464484
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_61
timestamp 1666464484
transform 1 0 6716 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_69
timestamp 1666464484
transform 1 0 7452 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_77
timestamp 1666464484
transform 1 0 8188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_81
timestamp 1666464484
transform 1 0 8556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1666464484
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_85
timestamp 1666464484
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_93
timestamp 1666464484
transform 1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_101
timestamp 1666464484
transform 1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_109
timestamp 1666464484
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_117
timestamp 1666464484
transform 1 0 11868 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_125
timestamp 1666464484
transform 1 0 12604 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_133
timestamp 1666464484
transform 1 0 13340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1666464484
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1666464484
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_141
timestamp 1666464484
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_149
timestamp 1666464484
transform 1 0 14812 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_157
timestamp 1666464484
transform 1 0 15548 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_165
timestamp 1666464484
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_173
timestamp 1666464484
transform 1 0 17020 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_181
timestamp 1666464484
transform 1 0 17756 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_189
timestamp 1666464484
transform 1 0 18492 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1666464484
transform 1 0 18860 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1666464484
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_197
timestamp 1666464484
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_205
timestamp 1666464484
transform 1 0 19964 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_213
timestamp 1666464484
transform 1 0 20700 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_221
timestamp 1666464484
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_229
timestamp 1666464484
transform 1 0 22172 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_237
timestamp 1666464484
transform 1 0 22908 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_245
timestamp 1666464484
transform 1 0 23644 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_249
timestamp 1666464484
transform 1 0 24012 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1666464484
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_253
timestamp 1666464484
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_261
timestamp 1666464484
transform 1 0 25116 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_269
timestamp 1666464484
transform 1 0 25852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_277
timestamp 1666464484
transform 1 0 26588 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_285
timestamp 1666464484
transform 1 0 27324 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_293
timestamp 1666464484
transform 1 0 28060 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_301
timestamp 1666464484
transform 1 0 28796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_305
timestamp 1666464484
transform 1 0 29164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1666464484
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_309
timestamp 1666464484
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_317
timestamp 1666464484
transform 1 0 30268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_325
timestamp 1666464484
transform 1 0 31004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_333
timestamp 1666464484
transform 1 0 31740 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_341
timestamp 1666464484
transform 1 0 32476 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_349
timestamp 1666464484
transform 1 0 33212 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_357
timestamp 1666464484
transform 1 0 33948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_361
timestamp 1666464484
transform 1 0 34316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1666464484
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_365
timestamp 1666464484
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_373
timestamp 1666464484
transform 1 0 35420 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_381
timestamp 1666464484
transform 1 0 36156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_389
timestamp 1666464484
transform 1 0 36892 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_397
timestamp 1666464484
transform 1 0 37628 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_405
timestamp 1666464484
transform 1 0 38364 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_413
timestamp 1666464484
transform 1 0 39100 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_417
timestamp 1666464484
transform 1 0 39468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1666464484
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_421
timestamp 1666464484
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_429
timestamp 1666464484
transform 1 0 40572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_437
timestamp 1666464484
transform 1 0 41308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_445
timestamp 1666464484
transform 1 0 42044 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_453
timestamp 1666464484
transform 1 0 42780 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_461
timestamp 1666464484
transform 1 0 43516 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_469
timestamp 1666464484
transform 1 0 44252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_473
timestamp 1666464484
transform 1 0 44620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1666464484
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_477
timestamp 1666464484
transform 1 0 44988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_485
timestamp 1666464484
transform 1 0 45724 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_493
timestamp 1666464484
transform 1 0 46460 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_501
timestamp 1666464484
transform 1 0 47196 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_509
timestamp 1666464484
transform 1 0 47932 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_517
timestamp 1666464484
transform 1 0 48668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_525
timestamp 1666464484
transform 1 0 49404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_529
timestamp 1666464484
transform 1 0 49772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1666464484
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_533
timestamp 1666464484
transform 1 0 50140 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_541
timestamp 1666464484
transform 1 0 50876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_549
timestamp 1666464484
transform 1 0 51612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_557
timestamp 1666464484
transform 1 0 52348 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_565
timestamp 1666464484
transform 1 0 53084 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_573
timestamp 1666464484
transform 1 0 53820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_581
timestamp 1666464484
transform 1 0 54556 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_585
timestamp 1666464484
transform 1 0 54924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1666464484
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_16_589
timestamp 1666464484
transform 1 0 55292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_597
timestamp 1666464484
transform 1 0 56028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_605
timestamp 1666464484
transform 1 0 56764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_16_613
timestamp 1666464484
transform 1 0 57500 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_16_621
timestamp 1666464484
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_17_3
timestamp 1666464484
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_11
timestamp 1666464484
transform 1 0 2116 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_19
timestamp 1666464484
transform 1 0 2852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_27
timestamp 1666464484
transform 1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_35
timestamp 1666464484
transform 1 0 4324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_43
timestamp 1666464484
transform 1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_51
timestamp 1666464484
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1666464484
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_57
timestamp 1666464484
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_65
timestamp 1666464484
transform 1 0 7084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_73
timestamp 1666464484
transform 1 0 7820 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_81
timestamp 1666464484
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_89
timestamp 1666464484
transform 1 0 9292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_97
timestamp 1666464484
transform 1 0 10028 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_105
timestamp 1666464484
transform 1 0 10764 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1666464484
transform 1 0 11132 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1666464484
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_113
timestamp 1666464484
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_121
timestamp 1666464484
transform 1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_129
timestamp 1666464484
transform 1 0 12972 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_137
timestamp 1666464484
transform 1 0 13708 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_145
timestamp 1666464484
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_153
timestamp 1666464484
transform 1 0 15180 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_161
timestamp 1666464484
transform 1 0 15916 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_165
timestamp 1666464484
transform 1 0 16284 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1666464484
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_169
timestamp 1666464484
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_177
timestamp 1666464484
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_185
timestamp 1666464484
transform 1 0 18124 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_193
timestamp 1666464484
transform 1 0 18860 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_201
timestamp 1666464484
transform 1 0 19596 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_209
timestamp 1666464484
transform 1 0 20332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_217
timestamp 1666464484
transform 1 0 21068 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1666464484
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1666464484
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_225
timestamp 1666464484
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_233
timestamp 1666464484
transform 1 0 22540 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_241
timestamp 1666464484
transform 1 0 23276 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_249
timestamp 1666464484
transform 1 0 24012 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_257
timestamp 1666464484
transform 1 0 24748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_265
timestamp 1666464484
transform 1 0 25484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_273
timestamp 1666464484
transform 1 0 26220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_277
timestamp 1666464484
transform 1 0 26588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1666464484
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_281
timestamp 1666464484
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_289
timestamp 1666464484
transform 1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_297
timestamp 1666464484
transform 1 0 28428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_305
timestamp 1666464484
transform 1 0 29164 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_313
timestamp 1666464484
transform 1 0 29900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_321
timestamp 1666464484
transform 1 0 30636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_329
timestamp 1666464484
transform 1 0 31372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_333
timestamp 1666464484
transform 1 0 31740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1666464484
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_337
timestamp 1666464484
transform 1 0 32108 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_345
timestamp 1666464484
transform 1 0 32844 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_353
timestamp 1666464484
transform 1 0 33580 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_361
timestamp 1666464484
transform 1 0 34316 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_369
timestamp 1666464484
transform 1 0 35052 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_377
timestamp 1666464484
transform 1 0 35788 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_385
timestamp 1666464484
transform 1 0 36524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_389
timestamp 1666464484
transform 1 0 36892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1666464484
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_393
timestamp 1666464484
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_401
timestamp 1666464484
transform 1 0 37996 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_409
timestamp 1666464484
transform 1 0 38732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_417
timestamp 1666464484
transform 1 0 39468 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_425
timestamp 1666464484
transform 1 0 40204 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_433
timestamp 1666464484
transform 1 0 40940 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_441
timestamp 1666464484
transform 1 0 41676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_445
timestamp 1666464484
transform 1 0 42044 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1666464484
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_449
timestamp 1666464484
transform 1 0 42412 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_457
timestamp 1666464484
transform 1 0 43148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_465
timestamp 1666464484
transform 1 0 43884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_473
timestamp 1666464484
transform 1 0 44620 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_481
timestamp 1666464484
transform 1 0 45356 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_489
timestamp 1666464484
transform 1 0 46092 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_497
timestamp 1666464484
transform 1 0 46828 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_501
timestamp 1666464484
transform 1 0 47196 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1666464484
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_505
timestamp 1666464484
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_513
timestamp 1666464484
transform 1 0 48300 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_521
timestamp 1666464484
transform 1 0 49036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_529
timestamp 1666464484
transform 1 0 49772 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_537
timestamp 1666464484
transform 1 0 50508 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_545
timestamp 1666464484
transform 1 0 51244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_553
timestamp 1666464484
transform 1 0 51980 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_557
timestamp 1666464484
transform 1 0 52348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1666464484
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_561
timestamp 1666464484
transform 1 0 52716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_569
timestamp 1666464484
transform 1 0 53452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_577
timestamp 1666464484
transform 1 0 54188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_585
timestamp 1666464484
transform 1 0 54924 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_593
timestamp 1666464484
transform 1 0 55660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_17_601
timestamp 1666464484
transform 1 0 56396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_609
timestamp 1666464484
transform 1 0 57132 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_613
timestamp 1666464484
transform 1 0 57500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1666464484
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_617
timestamp 1666464484
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_3
timestamp 1666464484
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_11
timestamp 1666464484
transform 1 0 2116 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_19
timestamp 1666464484
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1666464484
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_29
timestamp 1666464484
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_37
timestamp 1666464484
transform 1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_45
timestamp 1666464484
transform 1 0 5244 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_53
timestamp 1666464484
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_61
timestamp 1666464484
transform 1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_69
timestamp 1666464484
transform 1 0 7452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_77
timestamp 1666464484
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1666464484
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1666464484
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_85
timestamp 1666464484
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_93
timestamp 1666464484
transform 1 0 9660 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_101
timestamp 1666464484
transform 1 0 10396 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_109
timestamp 1666464484
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_117
timestamp 1666464484
transform 1 0 11868 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_125
timestamp 1666464484
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_133
timestamp 1666464484
transform 1 0 13340 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_137
timestamp 1666464484
transform 1 0 13708 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1666464484
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_141
timestamp 1666464484
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_149
timestamp 1666464484
transform 1 0 14812 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_157
timestamp 1666464484
transform 1 0 15548 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_165
timestamp 1666464484
transform 1 0 16284 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_173
timestamp 1666464484
transform 1 0 17020 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_181
timestamp 1666464484
transform 1 0 17756 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_189
timestamp 1666464484
transform 1 0 18492 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_193
timestamp 1666464484
transform 1 0 18860 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1666464484
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_197
timestamp 1666464484
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_205
timestamp 1666464484
transform 1 0 19964 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_213
timestamp 1666464484
transform 1 0 20700 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_221
timestamp 1666464484
transform 1 0 21436 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_229
timestamp 1666464484
transform 1 0 22172 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_237
timestamp 1666464484
transform 1 0 22908 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_245
timestamp 1666464484
transform 1 0 23644 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_249
timestamp 1666464484
transform 1 0 24012 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1666464484
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_253
timestamp 1666464484
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_261
timestamp 1666464484
transform 1 0 25116 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_269
timestamp 1666464484
transform 1 0 25852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_277
timestamp 1666464484
transform 1 0 26588 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_285
timestamp 1666464484
transform 1 0 27324 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_293
timestamp 1666464484
transform 1 0 28060 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_301
timestamp 1666464484
transform 1 0 28796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_305
timestamp 1666464484
transform 1 0 29164 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1666464484
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_309
timestamp 1666464484
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_317
timestamp 1666464484
transform 1 0 30268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_325
timestamp 1666464484
transform 1 0 31004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_333
timestamp 1666464484
transform 1 0 31740 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_341
timestamp 1666464484
transform 1 0 32476 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_349
timestamp 1666464484
transform 1 0 33212 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_357
timestamp 1666464484
transform 1 0 33948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_361
timestamp 1666464484
transform 1 0 34316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1666464484
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_365
timestamp 1666464484
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_373
timestamp 1666464484
transform 1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_381
timestamp 1666464484
transform 1 0 36156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_389
timestamp 1666464484
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_397
timestamp 1666464484
transform 1 0 37628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_405
timestamp 1666464484
transform 1 0 38364 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_413
timestamp 1666464484
transform 1 0 39100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_417
timestamp 1666464484
transform 1 0 39468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1666464484
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_421
timestamp 1666464484
transform 1 0 39836 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_429
timestamp 1666464484
transform 1 0 40572 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_437
timestamp 1666464484
transform 1 0 41308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_445
timestamp 1666464484
transform 1 0 42044 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_453
timestamp 1666464484
transform 1 0 42780 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_461
timestamp 1666464484
transform 1 0 43516 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_469
timestamp 1666464484
transform 1 0 44252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_473
timestamp 1666464484
transform 1 0 44620 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1666464484
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_477
timestamp 1666464484
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_485
timestamp 1666464484
transform 1 0 45724 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_493
timestamp 1666464484
transform 1 0 46460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_501
timestamp 1666464484
transform 1 0 47196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_509
timestamp 1666464484
transform 1 0 47932 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_517
timestamp 1666464484
transform 1 0 48668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_525
timestamp 1666464484
transform 1 0 49404 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_529
timestamp 1666464484
transform 1 0 49772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1666464484
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_533
timestamp 1666464484
transform 1 0 50140 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_541
timestamp 1666464484
transform 1 0 50876 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_549
timestamp 1666464484
transform 1 0 51612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_557
timestamp 1666464484
transform 1 0 52348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_565
timestamp 1666464484
transform 1 0 53084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_573
timestamp 1666464484
transform 1 0 53820 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_581
timestamp 1666464484
transform 1 0 54556 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_585
timestamp 1666464484
transform 1 0 54924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1666464484
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_589
timestamp 1666464484
transform 1 0 55292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_597
timestamp 1666464484
transform 1 0 56028 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_605
timestamp 1666464484
transform 1 0 56764 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_18_613
timestamp 1666464484
transform 1 0 57500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_18_621
timestamp 1666464484
transform 1 0 58236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_19_3
timestamp 1666464484
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_11
timestamp 1666464484
transform 1 0 2116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_19
timestamp 1666464484
transform 1 0 2852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_27
timestamp 1666464484
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_35
timestamp 1666464484
transform 1 0 4324 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_43
timestamp 1666464484
transform 1 0 5060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_51
timestamp 1666464484
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1666464484
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_57
timestamp 1666464484
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_65
timestamp 1666464484
transform 1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_73
timestamp 1666464484
transform 1 0 7820 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_81
timestamp 1666464484
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_89
timestamp 1666464484
transform 1 0 9292 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_97
timestamp 1666464484
transform 1 0 10028 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_105
timestamp 1666464484
transform 1 0 10764 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_109
timestamp 1666464484
transform 1 0 11132 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1666464484
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_113
timestamp 1666464484
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_121
timestamp 1666464484
transform 1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_129
timestamp 1666464484
transform 1 0 12972 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_137
timestamp 1666464484
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_145
timestamp 1666464484
transform 1 0 14444 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_153
timestamp 1666464484
transform 1 0 15180 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_161
timestamp 1666464484
transform 1 0 15916 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_165
timestamp 1666464484
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1666464484
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_169
timestamp 1666464484
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_177
timestamp 1666464484
transform 1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_185
timestamp 1666464484
transform 1 0 18124 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_193
timestamp 1666464484
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_201
timestamp 1666464484
transform 1 0 19596 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_209
timestamp 1666464484
transform 1 0 20332 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_217
timestamp 1666464484
transform 1 0 21068 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1666464484
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1666464484
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_225
timestamp 1666464484
transform 1 0 21804 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_233
timestamp 1666464484
transform 1 0 22540 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_241
timestamp 1666464484
transform 1 0 23276 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_249
timestamp 1666464484
transform 1 0 24012 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_257
timestamp 1666464484
transform 1 0 24748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_265
timestamp 1666464484
transform 1 0 25484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_273
timestamp 1666464484
transform 1 0 26220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_277
timestamp 1666464484
transform 1 0 26588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1666464484
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_281
timestamp 1666464484
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_289
timestamp 1666464484
transform 1 0 27692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_297
timestamp 1666464484
transform 1 0 28428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_305
timestamp 1666464484
transform 1 0 29164 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_313
timestamp 1666464484
transform 1 0 29900 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_321
timestamp 1666464484
transform 1 0 30636 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_329
timestamp 1666464484
transform 1 0 31372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_333
timestamp 1666464484
transform 1 0 31740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1666464484
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_337
timestamp 1666464484
transform 1 0 32108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_345
timestamp 1666464484
transform 1 0 32844 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_353
timestamp 1666464484
transform 1 0 33580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_361
timestamp 1666464484
transform 1 0 34316 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_369
timestamp 1666464484
transform 1 0 35052 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_377
timestamp 1666464484
transform 1 0 35788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_385
timestamp 1666464484
transform 1 0 36524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_389
timestamp 1666464484
transform 1 0 36892 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1666464484
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_393
timestamp 1666464484
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_401
timestamp 1666464484
transform 1 0 37996 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_409
timestamp 1666464484
transform 1 0 38732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_417
timestamp 1666464484
transform 1 0 39468 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_425
timestamp 1666464484
transform 1 0 40204 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_433
timestamp 1666464484
transform 1 0 40940 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_441
timestamp 1666464484
transform 1 0 41676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_445
timestamp 1666464484
transform 1 0 42044 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1666464484
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_449
timestamp 1666464484
transform 1 0 42412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_457
timestamp 1666464484
transform 1 0 43148 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_465
timestamp 1666464484
transform 1 0 43884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_473
timestamp 1666464484
transform 1 0 44620 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_481
timestamp 1666464484
transform 1 0 45356 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_489
timestamp 1666464484
transform 1 0 46092 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_497
timestamp 1666464484
transform 1 0 46828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_501
timestamp 1666464484
transform 1 0 47196 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1666464484
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_505
timestamp 1666464484
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_513
timestamp 1666464484
transform 1 0 48300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_521
timestamp 1666464484
transform 1 0 49036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_529
timestamp 1666464484
transform 1 0 49772 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_537
timestamp 1666464484
transform 1 0 50508 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_545
timestamp 1666464484
transform 1 0 51244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_553
timestamp 1666464484
transform 1 0 51980 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_557
timestamp 1666464484
transform 1 0 52348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1666464484
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_561
timestamp 1666464484
transform 1 0 52716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_569
timestamp 1666464484
transform 1 0 53452 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_577
timestamp 1666464484
transform 1 0 54188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_585
timestamp 1666464484
transform 1 0 54924 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_593
timestamp 1666464484
transform 1 0 55660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_19_601
timestamp 1666464484
transform 1 0 56396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_19_609
timestamp 1666464484
transform 1 0 57132 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_613
timestamp 1666464484
transform 1 0 57500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1666464484
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_617
timestamp 1666464484
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_3
timestamp 1666464484
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_11
timestamp 1666464484
transform 1 0 2116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_19
timestamp 1666464484
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1666464484
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_29
timestamp 1666464484
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_37
timestamp 1666464484
transform 1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_45
timestamp 1666464484
transform 1 0 5244 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_53
timestamp 1666464484
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_61
timestamp 1666464484
transform 1 0 6716 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_69
timestamp 1666464484
transform 1 0 7452 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_77
timestamp 1666464484
transform 1 0 8188 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1666464484
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1666464484
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_85
timestamp 1666464484
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_93
timestamp 1666464484
transform 1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_101
timestamp 1666464484
transform 1 0 10396 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_109
timestamp 1666464484
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_117
timestamp 1666464484
transform 1 0 11868 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_125
timestamp 1666464484
transform 1 0 12604 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_133
timestamp 1666464484
transform 1 0 13340 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_137
timestamp 1666464484
transform 1 0 13708 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1666464484
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_141
timestamp 1666464484
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_149
timestamp 1666464484
transform 1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_157
timestamp 1666464484
transform 1 0 15548 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_165
timestamp 1666464484
transform 1 0 16284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_173
timestamp 1666464484
transform 1 0 17020 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_181
timestamp 1666464484
transform 1 0 17756 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_189
timestamp 1666464484
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1666464484
transform 1 0 18860 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1666464484
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_197
timestamp 1666464484
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_205
timestamp 1666464484
transform 1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_213
timestamp 1666464484
transform 1 0 20700 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_221
timestamp 1666464484
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_229
timestamp 1666464484
transform 1 0 22172 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_237
timestamp 1666464484
transform 1 0 22908 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_245
timestamp 1666464484
transform 1 0 23644 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_249
timestamp 1666464484
transform 1 0 24012 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1666464484
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_253
timestamp 1666464484
transform 1 0 24380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_261
timestamp 1666464484
transform 1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_269
timestamp 1666464484
transform 1 0 25852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_277
timestamp 1666464484
transform 1 0 26588 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_285
timestamp 1666464484
transform 1 0 27324 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_293
timestamp 1666464484
transform 1 0 28060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_301
timestamp 1666464484
transform 1 0 28796 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_305
timestamp 1666464484
transform 1 0 29164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1666464484
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_309
timestamp 1666464484
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_317
timestamp 1666464484
transform 1 0 30268 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_325
timestamp 1666464484
transform 1 0 31004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_333
timestamp 1666464484
transform 1 0 31740 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_341
timestamp 1666464484
transform 1 0 32476 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_349
timestamp 1666464484
transform 1 0 33212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_357
timestamp 1666464484
transform 1 0 33948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_361
timestamp 1666464484
transform 1 0 34316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1666464484
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_365
timestamp 1666464484
transform 1 0 34684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_373
timestamp 1666464484
transform 1 0 35420 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_381
timestamp 1666464484
transform 1 0 36156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_389
timestamp 1666464484
transform 1 0 36892 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_397
timestamp 1666464484
transform 1 0 37628 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_405
timestamp 1666464484
transform 1 0 38364 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_413
timestamp 1666464484
transform 1 0 39100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_417
timestamp 1666464484
transform 1 0 39468 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1666464484
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_421
timestamp 1666464484
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_429
timestamp 1666464484
transform 1 0 40572 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_437
timestamp 1666464484
transform 1 0 41308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_445
timestamp 1666464484
transform 1 0 42044 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_453
timestamp 1666464484
transform 1 0 42780 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_461
timestamp 1666464484
transform 1 0 43516 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_469
timestamp 1666464484
transform 1 0 44252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_473
timestamp 1666464484
transform 1 0 44620 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1666464484
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_477
timestamp 1666464484
transform 1 0 44988 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_485
timestamp 1666464484
transform 1 0 45724 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_493
timestamp 1666464484
transform 1 0 46460 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_501
timestamp 1666464484
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_509
timestamp 1666464484
transform 1 0 47932 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_517
timestamp 1666464484
transform 1 0 48668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_525
timestamp 1666464484
transform 1 0 49404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_529
timestamp 1666464484
transform 1 0 49772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1666464484
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_533
timestamp 1666464484
transform 1 0 50140 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_541
timestamp 1666464484
transform 1 0 50876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_549
timestamp 1666464484
transform 1 0 51612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_557
timestamp 1666464484
transform 1 0 52348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_565
timestamp 1666464484
transform 1 0 53084 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_573
timestamp 1666464484
transform 1 0 53820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_581
timestamp 1666464484
transform 1 0 54556 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_585
timestamp 1666464484
transform 1 0 54924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1666464484
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_20_589
timestamp 1666464484
transform 1 0 55292 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_597
timestamp 1666464484
transform 1 0 56028 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_605
timestamp 1666464484
transform 1 0 56764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_613
timestamp 1666464484
transform 1 0 57500 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_621
timestamp 1666464484
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_21_3
timestamp 1666464484
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_11
timestamp 1666464484
transform 1 0 2116 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_19
timestamp 1666464484
transform 1 0 2852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_27
timestamp 1666464484
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_35
timestamp 1666464484
transform 1 0 4324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_43
timestamp 1666464484
transform 1 0 5060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_51
timestamp 1666464484
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1666464484
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_57
timestamp 1666464484
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_65
timestamp 1666464484
transform 1 0 7084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_73
timestamp 1666464484
transform 1 0 7820 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_81
timestamp 1666464484
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_89
timestamp 1666464484
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_97
timestamp 1666464484
transform 1 0 10028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_105
timestamp 1666464484
transform 1 0 10764 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1666464484
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1666464484
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_113
timestamp 1666464484
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_121
timestamp 1666464484
transform 1 0 12236 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_129
timestamp 1666464484
transform 1 0 12972 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_137
timestamp 1666464484
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_145
timestamp 1666464484
transform 1 0 14444 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_153
timestamp 1666464484
transform 1 0 15180 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_161
timestamp 1666464484
transform 1 0 15916 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_165
timestamp 1666464484
transform 1 0 16284 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1666464484
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_169
timestamp 1666464484
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_177
timestamp 1666464484
transform 1 0 17388 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_185
timestamp 1666464484
transform 1 0 18124 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_193
timestamp 1666464484
transform 1 0 18860 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_201
timestamp 1666464484
transform 1 0 19596 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_209
timestamp 1666464484
transform 1 0 20332 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_217
timestamp 1666464484
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1666464484
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1666464484
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_225
timestamp 1666464484
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_233
timestamp 1666464484
transform 1 0 22540 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_241
timestamp 1666464484
transform 1 0 23276 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_249
timestamp 1666464484
transform 1 0 24012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_257
timestamp 1666464484
transform 1 0 24748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_265
timestamp 1666464484
transform 1 0 25484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_273
timestamp 1666464484
transform 1 0 26220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_277
timestamp 1666464484
transform 1 0 26588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1666464484
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_281
timestamp 1666464484
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_289
timestamp 1666464484
transform 1 0 27692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_297
timestamp 1666464484
transform 1 0 28428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_305
timestamp 1666464484
transform 1 0 29164 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_313
timestamp 1666464484
transform 1 0 29900 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_321
timestamp 1666464484
transform 1 0 30636 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_329
timestamp 1666464484
transform 1 0 31372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_333
timestamp 1666464484
transform 1 0 31740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1666464484
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_337
timestamp 1666464484
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_345
timestamp 1666464484
transform 1 0 32844 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_353
timestamp 1666464484
transform 1 0 33580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_361
timestamp 1666464484
transform 1 0 34316 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_369
timestamp 1666464484
transform 1 0 35052 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_377
timestamp 1666464484
transform 1 0 35788 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_385
timestamp 1666464484
transform 1 0 36524 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_389
timestamp 1666464484
transform 1 0 36892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1666464484
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_393
timestamp 1666464484
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_401
timestamp 1666464484
transform 1 0 37996 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_409
timestamp 1666464484
transform 1 0 38732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_417
timestamp 1666464484
transform 1 0 39468 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_425
timestamp 1666464484
transform 1 0 40204 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_433
timestamp 1666464484
transform 1 0 40940 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_441
timestamp 1666464484
transform 1 0 41676 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_445
timestamp 1666464484
transform 1 0 42044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1666464484
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_449
timestamp 1666464484
transform 1 0 42412 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_457
timestamp 1666464484
transform 1 0 43148 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_465
timestamp 1666464484
transform 1 0 43884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_473
timestamp 1666464484
transform 1 0 44620 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_481
timestamp 1666464484
transform 1 0 45356 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_489
timestamp 1666464484
transform 1 0 46092 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_497
timestamp 1666464484
transform 1 0 46828 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_501
timestamp 1666464484
transform 1 0 47196 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1666464484
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_505
timestamp 1666464484
transform 1 0 47564 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_513
timestamp 1666464484
transform 1 0 48300 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_521
timestamp 1666464484
transform 1 0 49036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_529
timestamp 1666464484
transform 1 0 49772 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_537
timestamp 1666464484
transform 1 0 50508 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_545
timestamp 1666464484
transform 1 0 51244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_553
timestamp 1666464484
transform 1 0 51980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_557
timestamp 1666464484
transform 1 0 52348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1666464484
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_561
timestamp 1666464484
transform 1 0 52716 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_569
timestamp 1666464484
transform 1 0 53452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_577
timestamp 1666464484
transform 1 0 54188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_585
timestamp 1666464484
transform 1 0 54924 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_593
timestamp 1666464484
transform 1 0 55660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_21_601
timestamp 1666464484
transform 1 0 56396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_21_609
timestamp 1666464484
transform 1 0 57132 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_613
timestamp 1666464484
transform 1 0 57500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1666464484
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_617
timestamp 1666464484
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_3
timestamp 1666464484
transform 1 0 1380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_11
timestamp 1666464484
transform 1 0 2116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_19
timestamp 1666464484
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1666464484
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_29
timestamp 1666464484
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_37
timestamp 1666464484
transform 1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_45
timestamp 1666464484
transform 1 0 5244 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_53
timestamp 1666464484
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_61
timestamp 1666464484
transform 1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_69
timestamp 1666464484
transform 1 0 7452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_77
timestamp 1666464484
transform 1 0 8188 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_81
timestamp 1666464484
transform 1 0 8556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1666464484
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_85
timestamp 1666464484
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_93
timestamp 1666464484
transform 1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_101
timestamp 1666464484
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_109
timestamp 1666464484
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_117
timestamp 1666464484
transform 1 0 11868 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_125
timestamp 1666464484
transform 1 0 12604 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_133
timestamp 1666464484
transform 1 0 13340 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1666464484
transform 1 0 13708 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1666464484
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_141
timestamp 1666464484
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_149
timestamp 1666464484
transform 1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_157
timestamp 1666464484
transform 1 0 15548 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_165
timestamp 1666464484
transform 1 0 16284 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_173
timestamp 1666464484
transform 1 0 17020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_181
timestamp 1666464484
transform 1 0 17756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_189
timestamp 1666464484
transform 1 0 18492 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_193
timestamp 1666464484
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1666464484
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_197
timestamp 1666464484
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_205
timestamp 1666464484
transform 1 0 19964 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_213
timestamp 1666464484
transform 1 0 20700 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_221
timestamp 1666464484
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_229
timestamp 1666464484
transform 1 0 22172 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_237
timestamp 1666464484
transform 1 0 22908 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_245
timestamp 1666464484
transform 1 0 23644 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_249
timestamp 1666464484
transform 1 0 24012 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1666464484
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_253
timestamp 1666464484
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_261
timestamp 1666464484
transform 1 0 25116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_269
timestamp 1666464484
transform 1 0 25852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_277
timestamp 1666464484
transform 1 0 26588 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_285
timestamp 1666464484
transform 1 0 27324 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_293
timestamp 1666464484
transform 1 0 28060 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_301
timestamp 1666464484
transform 1 0 28796 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_305
timestamp 1666464484
transform 1 0 29164 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1666464484
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_309
timestamp 1666464484
transform 1 0 29532 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_317
timestamp 1666464484
transform 1 0 30268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_325
timestamp 1666464484
transform 1 0 31004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_333
timestamp 1666464484
transform 1 0 31740 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_341
timestamp 1666464484
transform 1 0 32476 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_349
timestamp 1666464484
transform 1 0 33212 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_357
timestamp 1666464484
transform 1 0 33948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_361
timestamp 1666464484
transform 1 0 34316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1666464484
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_365
timestamp 1666464484
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_373
timestamp 1666464484
transform 1 0 35420 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_381
timestamp 1666464484
transform 1 0 36156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_389
timestamp 1666464484
transform 1 0 36892 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_397
timestamp 1666464484
transform 1 0 37628 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_405
timestamp 1666464484
transform 1 0 38364 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_413
timestamp 1666464484
transform 1 0 39100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_417
timestamp 1666464484
transform 1 0 39468 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1666464484
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_421
timestamp 1666464484
transform 1 0 39836 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_429
timestamp 1666464484
transform 1 0 40572 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_437
timestamp 1666464484
transform 1 0 41308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_445
timestamp 1666464484
transform 1 0 42044 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_453
timestamp 1666464484
transform 1 0 42780 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_461
timestamp 1666464484
transform 1 0 43516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_469
timestamp 1666464484
transform 1 0 44252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_473
timestamp 1666464484
transform 1 0 44620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1666464484
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_477
timestamp 1666464484
transform 1 0 44988 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_485
timestamp 1666464484
transform 1 0 45724 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_493
timestamp 1666464484
transform 1 0 46460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_501
timestamp 1666464484
transform 1 0 47196 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_509
timestamp 1666464484
transform 1 0 47932 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_517
timestamp 1666464484
transform 1 0 48668 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_525
timestamp 1666464484
transform 1 0 49404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_529
timestamp 1666464484
transform 1 0 49772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1666464484
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_533
timestamp 1666464484
transform 1 0 50140 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_541
timestamp 1666464484
transform 1 0 50876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_549
timestamp 1666464484
transform 1 0 51612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_557
timestamp 1666464484
transform 1 0 52348 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_565
timestamp 1666464484
transform 1 0 53084 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_573
timestamp 1666464484
transform 1 0 53820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_581
timestamp 1666464484
transform 1 0 54556 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_585
timestamp 1666464484
transform 1 0 54924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1666464484
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_22_589
timestamp 1666464484
transform 1 0 55292 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_597
timestamp 1666464484
transform 1 0 56028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_605
timestamp 1666464484
transform 1 0 56764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_22_613
timestamp 1666464484
transform 1 0 57500 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_621
timestamp 1666464484
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_23_3
timestamp 1666464484
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_11
timestamp 1666464484
transform 1 0 2116 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_19
timestamp 1666464484
transform 1 0 2852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_27
timestamp 1666464484
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_35
timestamp 1666464484
transform 1 0 4324 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_43
timestamp 1666464484
transform 1 0 5060 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_51
timestamp 1666464484
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1666464484
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_57
timestamp 1666464484
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_65
timestamp 1666464484
transform 1 0 7084 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_73
timestamp 1666464484
transform 1 0 7820 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_81
timestamp 1666464484
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_89
timestamp 1666464484
transform 1 0 9292 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_97
timestamp 1666464484
transform 1 0 10028 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_105
timestamp 1666464484
transform 1 0 10764 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_109
timestamp 1666464484
transform 1 0 11132 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1666464484
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_113
timestamp 1666464484
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_121
timestamp 1666464484
transform 1 0 12236 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_129
timestamp 1666464484
transform 1 0 12972 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_137
timestamp 1666464484
transform 1 0 13708 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_145
timestamp 1666464484
transform 1 0 14444 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_153
timestamp 1666464484
transform 1 0 15180 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_161
timestamp 1666464484
transform 1 0 15916 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_165
timestamp 1666464484
transform 1 0 16284 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1666464484
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_169
timestamp 1666464484
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_177
timestamp 1666464484
transform 1 0 17388 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_185
timestamp 1666464484
transform 1 0 18124 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_193
timestamp 1666464484
transform 1 0 18860 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_201
timestamp 1666464484
transform 1 0 19596 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_209
timestamp 1666464484
transform 1 0 20332 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_217
timestamp 1666464484
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1666464484
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1666464484
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_225
timestamp 1666464484
transform 1 0 21804 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_233
timestamp 1666464484
transform 1 0 22540 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_241
timestamp 1666464484
transform 1 0 23276 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_249
timestamp 1666464484
transform 1 0 24012 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_257
timestamp 1666464484
transform 1 0 24748 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_265
timestamp 1666464484
transform 1 0 25484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_273
timestamp 1666464484
transform 1 0 26220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_277
timestamp 1666464484
transform 1 0 26588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1666464484
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_281
timestamp 1666464484
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_289
timestamp 1666464484
transform 1 0 27692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_297
timestamp 1666464484
transform 1 0 28428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_305
timestamp 1666464484
transform 1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_313
timestamp 1666464484
transform 1 0 29900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_321
timestamp 1666464484
transform 1 0 30636 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_329
timestamp 1666464484
transform 1 0 31372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_333
timestamp 1666464484
transform 1 0 31740 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1666464484
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_337
timestamp 1666464484
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_345
timestamp 1666464484
transform 1 0 32844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_353
timestamp 1666464484
transform 1 0 33580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_361
timestamp 1666464484
transform 1 0 34316 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_369
timestamp 1666464484
transform 1 0 35052 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_377
timestamp 1666464484
transform 1 0 35788 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_385
timestamp 1666464484
transform 1 0 36524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_389
timestamp 1666464484
transform 1 0 36892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1666464484
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_393
timestamp 1666464484
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_401
timestamp 1666464484
transform 1 0 37996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_409
timestamp 1666464484
transform 1 0 38732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_417
timestamp 1666464484
transform 1 0 39468 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_425
timestamp 1666464484
transform 1 0 40204 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_433
timestamp 1666464484
transform 1 0 40940 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_441
timestamp 1666464484
transform 1 0 41676 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_445
timestamp 1666464484
transform 1 0 42044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1666464484
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_449
timestamp 1666464484
transform 1 0 42412 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_457
timestamp 1666464484
transform 1 0 43148 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_465
timestamp 1666464484
transform 1 0 43884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_473
timestamp 1666464484
transform 1 0 44620 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_481
timestamp 1666464484
transform 1 0 45356 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_489
timestamp 1666464484
transform 1 0 46092 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_497
timestamp 1666464484
transform 1 0 46828 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_501
timestamp 1666464484
transform 1 0 47196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1666464484
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_505
timestamp 1666464484
transform 1 0 47564 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_513
timestamp 1666464484
transform 1 0 48300 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_521
timestamp 1666464484
transform 1 0 49036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_529
timestamp 1666464484
transform 1 0 49772 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_537
timestamp 1666464484
transform 1 0 50508 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_545
timestamp 1666464484
transform 1 0 51244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_553
timestamp 1666464484
transform 1 0 51980 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_557
timestamp 1666464484
transform 1 0 52348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1666464484
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_561
timestamp 1666464484
transform 1 0 52716 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_569
timestamp 1666464484
transform 1 0 53452 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_577
timestamp 1666464484
transform 1 0 54188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_585
timestamp 1666464484
transform 1 0 54924 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_593
timestamp 1666464484
transform 1 0 55660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_23_601
timestamp 1666464484
transform 1 0 56396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_23_609
timestamp 1666464484
transform 1 0 57132 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_613
timestamp 1666464484
transform 1 0 57500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1666464484
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_617
timestamp 1666464484
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_3
timestamp 1666464484
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_11
timestamp 1666464484
transform 1 0 2116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_19
timestamp 1666464484
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1666464484
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_29
timestamp 1666464484
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_37
timestamp 1666464484
transform 1 0 4508 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_45
timestamp 1666464484
transform 1 0 5244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_53
timestamp 1666464484
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_61
timestamp 1666464484
transform 1 0 6716 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_69
timestamp 1666464484
transform 1 0 7452 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_77
timestamp 1666464484
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_81
timestamp 1666464484
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1666464484
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_85
timestamp 1666464484
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_93
timestamp 1666464484
transform 1 0 9660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_101
timestamp 1666464484
transform 1 0 10396 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_109
timestamp 1666464484
transform 1 0 11132 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_117
timestamp 1666464484
transform 1 0 11868 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_125
timestamp 1666464484
transform 1 0 12604 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_133
timestamp 1666464484
transform 1 0 13340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_137
timestamp 1666464484
transform 1 0 13708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1666464484
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_141
timestamp 1666464484
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_149
timestamp 1666464484
transform 1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_157
timestamp 1666464484
transform 1 0 15548 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_165
timestamp 1666464484
transform 1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_173
timestamp 1666464484
transform 1 0 17020 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_181
timestamp 1666464484
transform 1 0 17756 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_189
timestamp 1666464484
transform 1 0 18492 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1666464484
transform 1 0 18860 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1666464484
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_197
timestamp 1666464484
transform 1 0 19228 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_205
timestamp 1666464484
transform 1 0 19964 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_213
timestamp 1666464484
transform 1 0 20700 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_221
timestamp 1666464484
transform 1 0 21436 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_229
timestamp 1666464484
transform 1 0 22172 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_237
timestamp 1666464484
transform 1 0 22908 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_245
timestamp 1666464484
transform 1 0 23644 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_249
timestamp 1666464484
transform 1 0 24012 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1666464484
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_253
timestamp 1666464484
transform 1 0 24380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_261
timestamp 1666464484
transform 1 0 25116 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_269
timestamp 1666464484
transform 1 0 25852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_277
timestamp 1666464484
transform 1 0 26588 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_285
timestamp 1666464484
transform 1 0 27324 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_293
timestamp 1666464484
transform 1 0 28060 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_301
timestamp 1666464484
transform 1 0 28796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_305
timestamp 1666464484
transform 1 0 29164 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1666464484
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_309
timestamp 1666464484
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_317
timestamp 1666464484
transform 1 0 30268 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_325
timestamp 1666464484
transform 1 0 31004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_333
timestamp 1666464484
transform 1 0 31740 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_341
timestamp 1666464484
transform 1 0 32476 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_349
timestamp 1666464484
transform 1 0 33212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_357
timestamp 1666464484
transform 1 0 33948 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_361
timestamp 1666464484
transform 1 0 34316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1666464484
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_365
timestamp 1666464484
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_373
timestamp 1666464484
transform 1 0 35420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_381
timestamp 1666464484
transform 1 0 36156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_389
timestamp 1666464484
transform 1 0 36892 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_397
timestamp 1666464484
transform 1 0 37628 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_405
timestamp 1666464484
transform 1 0 38364 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_413
timestamp 1666464484
transform 1 0 39100 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_417
timestamp 1666464484
transform 1 0 39468 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1666464484
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_421
timestamp 1666464484
transform 1 0 39836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_429
timestamp 1666464484
transform 1 0 40572 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_437
timestamp 1666464484
transform 1 0 41308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_445
timestamp 1666464484
transform 1 0 42044 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_453
timestamp 1666464484
transform 1 0 42780 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_461
timestamp 1666464484
transform 1 0 43516 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_469
timestamp 1666464484
transform 1 0 44252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_473
timestamp 1666464484
transform 1 0 44620 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1666464484
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_477
timestamp 1666464484
transform 1 0 44988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_485
timestamp 1666464484
transform 1 0 45724 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_493
timestamp 1666464484
transform 1 0 46460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_501
timestamp 1666464484
transform 1 0 47196 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_509
timestamp 1666464484
transform 1 0 47932 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_517
timestamp 1666464484
transform 1 0 48668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_525
timestamp 1666464484
transform 1 0 49404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_529
timestamp 1666464484
transform 1 0 49772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1666464484
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_533
timestamp 1666464484
transform 1 0 50140 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_541
timestamp 1666464484
transform 1 0 50876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_549
timestamp 1666464484
transform 1 0 51612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_557
timestamp 1666464484
transform 1 0 52348 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_565
timestamp 1666464484
transform 1 0 53084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_573
timestamp 1666464484
transform 1 0 53820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_581
timestamp 1666464484
transform 1 0 54556 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_585
timestamp 1666464484
transform 1 0 54924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1666464484
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_24_589
timestamp 1666464484
transform 1 0 55292 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_597
timestamp 1666464484
transform 1 0 56028 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_605
timestamp 1666464484
transform 1 0 56764 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_24_613
timestamp 1666464484
transform 1 0 57500 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_621
timestamp 1666464484
transform 1 0 58236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_25_3
timestamp 1666464484
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_11
timestamp 1666464484
transform 1 0 2116 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_19
timestamp 1666464484
transform 1 0 2852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_27
timestamp 1666464484
transform 1 0 3588 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_35
timestamp 1666464484
transform 1 0 4324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_43
timestamp 1666464484
transform 1 0 5060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_51
timestamp 1666464484
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1666464484
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_57
timestamp 1666464484
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_65
timestamp 1666464484
transform 1 0 7084 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_73
timestamp 1666464484
transform 1 0 7820 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_81
timestamp 1666464484
transform 1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_89
timestamp 1666464484
transform 1 0 9292 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_97
timestamp 1666464484
transform 1 0 10028 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_105
timestamp 1666464484
transform 1 0 10764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_109
timestamp 1666464484
transform 1 0 11132 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1666464484
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_113
timestamp 1666464484
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_121
timestamp 1666464484
transform 1 0 12236 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_129
timestamp 1666464484
transform 1 0 12972 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_137
timestamp 1666464484
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_145
timestamp 1666464484
transform 1 0 14444 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_153
timestamp 1666464484
transform 1 0 15180 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_161
timestamp 1666464484
transform 1 0 15916 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_165
timestamp 1666464484
transform 1 0 16284 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1666464484
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_169
timestamp 1666464484
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_177
timestamp 1666464484
transform 1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_185
timestamp 1666464484
transform 1 0 18124 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_193
timestamp 1666464484
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_201
timestamp 1666464484
transform 1 0 19596 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_209
timestamp 1666464484
transform 1 0 20332 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_217
timestamp 1666464484
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1666464484
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1666464484
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_225
timestamp 1666464484
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_233
timestamp 1666464484
transform 1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_241
timestamp 1666464484
transform 1 0 23276 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_249
timestamp 1666464484
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_257
timestamp 1666464484
transform 1 0 24748 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_265
timestamp 1666464484
transform 1 0 25484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_273
timestamp 1666464484
transform 1 0 26220 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_277
timestamp 1666464484
transform 1 0 26588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1666464484
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_281
timestamp 1666464484
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_289
timestamp 1666464484
transform 1 0 27692 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_297
timestamp 1666464484
transform 1 0 28428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_305
timestamp 1666464484
transform 1 0 29164 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_313
timestamp 1666464484
transform 1 0 29900 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_321
timestamp 1666464484
transform 1 0 30636 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_329
timestamp 1666464484
transform 1 0 31372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_333
timestamp 1666464484
transform 1 0 31740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1666464484
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_337
timestamp 1666464484
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_345
timestamp 1666464484
transform 1 0 32844 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_353
timestamp 1666464484
transform 1 0 33580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_361
timestamp 1666464484
transform 1 0 34316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_369
timestamp 1666464484
transform 1 0 35052 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_377
timestamp 1666464484
transform 1 0 35788 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_385
timestamp 1666464484
transform 1 0 36524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_389
timestamp 1666464484
transform 1 0 36892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1666464484
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_393
timestamp 1666464484
transform 1 0 37260 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_401
timestamp 1666464484
transform 1 0 37996 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_409
timestamp 1666464484
transform 1 0 38732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_417
timestamp 1666464484
transform 1 0 39468 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_425
timestamp 1666464484
transform 1 0 40204 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_433
timestamp 1666464484
transform 1 0 40940 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_441
timestamp 1666464484
transform 1 0 41676 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_445
timestamp 1666464484
transform 1 0 42044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1666464484
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_449
timestamp 1666464484
transform 1 0 42412 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_457
timestamp 1666464484
transform 1 0 43148 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_465
timestamp 1666464484
transform 1 0 43884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_473
timestamp 1666464484
transform 1 0 44620 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_481
timestamp 1666464484
transform 1 0 45356 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_489
timestamp 1666464484
transform 1 0 46092 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_497
timestamp 1666464484
transform 1 0 46828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_501
timestamp 1666464484
transform 1 0 47196 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1666464484
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_505
timestamp 1666464484
transform 1 0 47564 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_513
timestamp 1666464484
transform 1 0 48300 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_521
timestamp 1666464484
transform 1 0 49036 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_529
timestamp 1666464484
transform 1 0 49772 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_537
timestamp 1666464484
transform 1 0 50508 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_545
timestamp 1666464484
transform 1 0 51244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_553
timestamp 1666464484
transform 1 0 51980 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_557
timestamp 1666464484
transform 1 0 52348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1666464484
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_561
timestamp 1666464484
transform 1 0 52716 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_569
timestamp 1666464484
transform 1 0 53452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_577
timestamp 1666464484
transform 1 0 54188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_585
timestamp 1666464484
transform 1 0 54924 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_593
timestamp 1666464484
transform 1 0 55660 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_25_601
timestamp 1666464484
transform 1 0 56396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_609
timestamp 1666464484
transform 1 0 57132 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_613
timestamp 1666464484
transform 1 0 57500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1666464484
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_617
timestamp 1666464484
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_3
timestamp 1666464484
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_11
timestamp 1666464484
transform 1 0 2116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_19
timestamp 1666464484
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1666464484
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_29
timestamp 1666464484
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_37
timestamp 1666464484
transform 1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_45
timestamp 1666464484
transform 1 0 5244 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_53
timestamp 1666464484
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_61
timestamp 1666464484
transform 1 0 6716 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_69
timestamp 1666464484
transform 1 0 7452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_77
timestamp 1666464484
transform 1 0 8188 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_81
timestamp 1666464484
transform 1 0 8556 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1666464484
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_85
timestamp 1666464484
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_93
timestamp 1666464484
transform 1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_101
timestamp 1666464484
transform 1 0 10396 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_109
timestamp 1666464484
transform 1 0 11132 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_117
timestamp 1666464484
transform 1 0 11868 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_125
timestamp 1666464484
transform 1 0 12604 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_133
timestamp 1666464484
transform 1 0 13340 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_137
timestamp 1666464484
transform 1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1666464484
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_141
timestamp 1666464484
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_149
timestamp 1666464484
transform 1 0 14812 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_157
timestamp 1666464484
transform 1 0 15548 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_165
timestamp 1666464484
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_173
timestamp 1666464484
transform 1 0 17020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_181
timestamp 1666464484
transform 1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_189
timestamp 1666464484
transform 1 0 18492 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_193
timestamp 1666464484
transform 1 0 18860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1666464484
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_197
timestamp 1666464484
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_205
timestamp 1666464484
transform 1 0 19964 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_213
timestamp 1666464484
transform 1 0 20700 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_221
timestamp 1666464484
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_229
timestamp 1666464484
transform 1 0 22172 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_237
timestamp 1666464484
transform 1 0 22908 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_245
timestamp 1666464484
transform 1 0 23644 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_249
timestamp 1666464484
transform 1 0 24012 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1666464484
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_253
timestamp 1666464484
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_261
timestamp 1666464484
transform 1 0 25116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_269
timestamp 1666464484
transform 1 0 25852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_277
timestamp 1666464484
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_285
timestamp 1666464484
transform 1 0 27324 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_293
timestamp 1666464484
transform 1 0 28060 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_301
timestamp 1666464484
transform 1 0 28796 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_305
timestamp 1666464484
transform 1 0 29164 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1666464484
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_309
timestamp 1666464484
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_317
timestamp 1666464484
transform 1 0 30268 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_325
timestamp 1666464484
transform 1 0 31004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_333
timestamp 1666464484
transform 1 0 31740 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_341
timestamp 1666464484
transform 1 0 32476 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_349
timestamp 1666464484
transform 1 0 33212 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_357
timestamp 1666464484
transform 1 0 33948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_361
timestamp 1666464484
transform 1 0 34316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1666464484
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_365
timestamp 1666464484
transform 1 0 34684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_373
timestamp 1666464484
transform 1 0 35420 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_381
timestamp 1666464484
transform 1 0 36156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_389
timestamp 1666464484
transform 1 0 36892 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_397
timestamp 1666464484
transform 1 0 37628 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_405
timestamp 1666464484
transform 1 0 38364 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_413
timestamp 1666464484
transform 1 0 39100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_417
timestamp 1666464484
transform 1 0 39468 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1666464484
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_421
timestamp 1666464484
transform 1 0 39836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_429
timestamp 1666464484
transform 1 0 40572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_437
timestamp 1666464484
transform 1 0 41308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_445
timestamp 1666464484
transform 1 0 42044 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_453
timestamp 1666464484
transform 1 0 42780 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_461
timestamp 1666464484
transform 1 0 43516 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_469
timestamp 1666464484
transform 1 0 44252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_473
timestamp 1666464484
transform 1 0 44620 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1666464484
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_477
timestamp 1666464484
transform 1 0 44988 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_485
timestamp 1666464484
transform 1 0 45724 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_493
timestamp 1666464484
transform 1 0 46460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_501
timestamp 1666464484
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_509
timestamp 1666464484
transform 1 0 47932 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_517
timestamp 1666464484
transform 1 0 48668 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_525
timestamp 1666464484
transform 1 0 49404 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_529
timestamp 1666464484
transform 1 0 49772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1666464484
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_533
timestamp 1666464484
transform 1 0 50140 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_541
timestamp 1666464484
transform 1 0 50876 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_549
timestamp 1666464484
transform 1 0 51612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_557
timestamp 1666464484
transform 1 0 52348 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_565
timestamp 1666464484
transform 1 0 53084 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_573
timestamp 1666464484
transform 1 0 53820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_581
timestamp 1666464484
transform 1 0 54556 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_585
timestamp 1666464484
transform 1 0 54924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1666464484
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_26_589
timestamp 1666464484
transform 1 0 55292 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_597
timestamp 1666464484
transform 1 0 56028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_605
timestamp 1666464484
transform 1 0 56764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_26_613
timestamp 1666464484
transform 1 0 57500 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_621
timestamp 1666464484
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_27_3
timestamp 1666464484
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_11
timestamp 1666464484
transform 1 0 2116 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_19
timestamp 1666464484
transform 1 0 2852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_27
timestamp 1666464484
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_35
timestamp 1666464484
transform 1 0 4324 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_43
timestamp 1666464484
transform 1 0 5060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_51
timestamp 1666464484
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1666464484
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_57
timestamp 1666464484
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_65
timestamp 1666464484
transform 1 0 7084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_73
timestamp 1666464484
transform 1 0 7820 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_81
timestamp 1666464484
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_89
timestamp 1666464484
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_97
timestamp 1666464484
transform 1 0 10028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_105
timestamp 1666464484
transform 1 0 10764 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1666464484
transform 1 0 11132 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1666464484
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_113
timestamp 1666464484
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_121
timestamp 1666464484
transform 1 0 12236 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_129
timestamp 1666464484
transform 1 0 12972 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_137
timestamp 1666464484
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_145
timestamp 1666464484
transform 1 0 14444 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_153
timestamp 1666464484
transform 1 0 15180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_161
timestamp 1666464484
transform 1 0 15916 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1666464484
transform 1 0 16284 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1666464484
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_169
timestamp 1666464484
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_177
timestamp 1666464484
transform 1 0 17388 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_185
timestamp 1666464484
transform 1 0 18124 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_193
timestamp 1666464484
transform 1 0 18860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_201
timestamp 1666464484
transform 1 0 19596 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_209
timestamp 1666464484
transform 1 0 20332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_217
timestamp 1666464484
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1666464484
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1666464484
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_225
timestamp 1666464484
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_233
timestamp 1666464484
transform 1 0 22540 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_241
timestamp 1666464484
transform 1 0 23276 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_249
timestamp 1666464484
transform 1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_257
timestamp 1666464484
transform 1 0 24748 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_265
timestamp 1666464484
transform 1 0 25484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_273
timestamp 1666464484
transform 1 0 26220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_277
timestamp 1666464484
transform 1 0 26588 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1666464484
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_281
timestamp 1666464484
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_289
timestamp 1666464484
transform 1 0 27692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_297
timestamp 1666464484
transform 1 0 28428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_305
timestamp 1666464484
transform 1 0 29164 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_313
timestamp 1666464484
transform 1 0 29900 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_321
timestamp 1666464484
transform 1 0 30636 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_329
timestamp 1666464484
transform 1 0 31372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_333
timestamp 1666464484
transform 1 0 31740 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1666464484
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_337
timestamp 1666464484
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_345
timestamp 1666464484
transform 1 0 32844 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_353
timestamp 1666464484
transform 1 0 33580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_361
timestamp 1666464484
transform 1 0 34316 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_369
timestamp 1666464484
transform 1 0 35052 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_377
timestamp 1666464484
transform 1 0 35788 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_385
timestamp 1666464484
transform 1 0 36524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_389
timestamp 1666464484
transform 1 0 36892 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1666464484
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_393
timestamp 1666464484
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_401
timestamp 1666464484
transform 1 0 37996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_409
timestamp 1666464484
transform 1 0 38732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_417
timestamp 1666464484
transform 1 0 39468 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_425
timestamp 1666464484
transform 1 0 40204 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_433
timestamp 1666464484
transform 1 0 40940 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_441
timestamp 1666464484
transform 1 0 41676 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_445
timestamp 1666464484
transform 1 0 42044 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1666464484
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_449
timestamp 1666464484
transform 1 0 42412 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_457
timestamp 1666464484
transform 1 0 43148 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_465
timestamp 1666464484
transform 1 0 43884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_473
timestamp 1666464484
transform 1 0 44620 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_481
timestamp 1666464484
transform 1 0 45356 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_489
timestamp 1666464484
transform 1 0 46092 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_497
timestamp 1666464484
transform 1 0 46828 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_501
timestamp 1666464484
transform 1 0 47196 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1666464484
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_505
timestamp 1666464484
transform 1 0 47564 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_513
timestamp 1666464484
transform 1 0 48300 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_521
timestamp 1666464484
transform 1 0 49036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_529
timestamp 1666464484
transform 1 0 49772 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_537
timestamp 1666464484
transform 1 0 50508 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_545
timestamp 1666464484
transform 1 0 51244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_553
timestamp 1666464484
transform 1 0 51980 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_557
timestamp 1666464484
transform 1 0 52348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1666464484
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_561
timestamp 1666464484
transform 1 0 52716 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_569
timestamp 1666464484
transform 1 0 53452 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_577
timestamp 1666464484
transform 1 0 54188 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_585
timestamp 1666464484
transform 1 0 54924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_593
timestamp 1666464484
transform 1 0 55660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_601
timestamp 1666464484
transform 1 0 56396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_27_609
timestamp 1666464484
transform 1 0 57132 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_613
timestamp 1666464484
transform 1 0 57500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1666464484
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_617
timestamp 1666464484
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_3
timestamp 1666464484
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_11
timestamp 1666464484
transform 1 0 2116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_19
timestamp 1666464484
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1666464484
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_29
timestamp 1666464484
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_37
timestamp 1666464484
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_45
timestamp 1666464484
transform 1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_53
timestamp 1666464484
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_61
timestamp 1666464484
transform 1 0 6716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_69
timestamp 1666464484
transform 1 0 7452 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_77
timestamp 1666464484
transform 1 0 8188 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_81
timestamp 1666464484
transform 1 0 8556 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1666464484
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_85
timestamp 1666464484
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_93
timestamp 1666464484
transform 1 0 9660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_101
timestamp 1666464484
transform 1 0 10396 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_109
timestamp 1666464484
transform 1 0 11132 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_117
timestamp 1666464484
transform 1 0 11868 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_125
timestamp 1666464484
transform 1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_133
timestamp 1666464484
transform 1 0 13340 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_137
timestamp 1666464484
transform 1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1666464484
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_141
timestamp 1666464484
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_149
timestamp 1666464484
transform 1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_157
timestamp 1666464484
transform 1 0 15548 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_165
timestamp 1666464484
transform 1 0 16284 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_173
timestamp 1666464484
transform 1 0 17020 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_181
timestamp 1666464484
transform 1 0 17756 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_189
timestamp 1666464484
transform 1 0 18492 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1666464484
transform 1 0 18860 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1666464484
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_197
timestamp 1666464484
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_205
timestamp 1666464484
transform 1 0 19964 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_213
timestamp 1666464484
transform 1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_221
timestamp 1666464484
transform 1 0 21436 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_229
timestamp 1666464484
transform 1 0 22172 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_237
timestamp 1666464484
transform 1 0 22908 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_245
timestamp 1666464484
transform 1 0 23644 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_249
timestamp 1666464484
transform 1 0 24012 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1666464484
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_253
timestamp 1666464484
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_261
timestamp 1666464484
transform 1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_269
timestamp 1666464484
transform 1 0 25852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_277
timestamp 1666464484
transform 1 0 26588 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_285
timestamp 1666464484
transform 1 0 27324 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_293
timestamp 1666464484
transform 1 0 28060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_301
timestamp 1666464484
transform 1 0 28796 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_305
timestamp 1666464484
transform 1 0 29164 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1666464484
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_309
timestamp 1666464484
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_317
timestamp 1666464484
transform 1 0 30268 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_325
timestamp 1666464484
transform 1 0 31004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_333
timestamp 1666464484
transform 1 0 31740 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_341
timestamp 1666464484
transform 1 0 32476 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_349
timestamp 1666464484
transform 1 0 33212 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_357
timestamp 1666464484
transform 1 0 33948 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_361
timestamp 1666464484
transform 1 0 34316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1666464484
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_365
timestamp 1666464484
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_373
timestamp 1666464484
transform 1 0 35420 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_381
timestamp 1666464484
transform 1 0 36156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_389
timestamp 1666464484
transform 1 0 36892 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_397
timestamp 1666464484
transform 1 0 37628 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_405
timestamp 1666464484
transform 1 0 38364 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_413
timestamp 1666464484
transform 1 0 39100 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_417
timestamp 1666464484
transform 1 0 39468 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1666464484
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_421
timestamp 1666464484
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_429
timestamp 1666464484
transform 1 0 40572 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_437
timestamp 1666464484
transform 1 0 41308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_445
timestamp 1666464484
transform 1 0 42044 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_453
timestamp 1666464484
transform 1 0 42780 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_461
timestamp 1666464484
transform 1 0 43516 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_469
timestamp 1666464484
transform 1 0 44252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_473
timestamp 1666464484
transform 1 0 44620 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1666464484
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_477
timestamp 1666464484
transform 1 0 44988 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_485
timestamp 1666464484
transform 1 0 45724 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_493
timestamp 1666464484
transform 1 0 46460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_501
timestamp 1666464484
transform 1 0 47196 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_509
timestamp 1666464484
transform 1 0 47932 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_517
timestamp 1666464484
transform 1 0 48668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_525
timestamp 1666464484
transform 1 0 49404 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_529
timestamp 1666464484
transform 1 0 49772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1666464484
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_533
timestamp 1666464484
transform 1 0 50140 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_541
timestamp 1666464484
transform 1 0 50876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_549
timestamp 1666464484
transform 1 0 51612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_557
timestamp 1666464484
transform 1 0 52348 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_565
timestamp 1666464484
transform 1 0 53084 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_573
timestamp 1666464484
transform 1 0 53820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_581
timestamp 1666464484
transform 1 0 54556 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_585
timestamp 1666464484
transform 1 0 54924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1666464484
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_589
timestamp 1666464484
transform 1 0 55292 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_597
timestamp 1666464484
transform 1 0 56028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_605
timestamp 1666464484
transform 1 0 56764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_28_613
timestamp 1666464484
transform 1 0 57500 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_28_621
timestamp 1666464484
transform 1 0 58236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_29_3
timestamp 1666464484
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_11
timestamp 1666464484
transform 1 0 2116 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_19
timestamp 1666464484
transform 1 0 2852 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_27
timestamp 1666464484
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_35
timestamp 1666464484
transform 1 0 4324 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_43
timestamp 1666464484
transform 1 0 5060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_51
timestamp 1666464484
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1666464484
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_57
timestamp 1666464484
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_65
timestamp 1666464484
transform 1 0 7084 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_73
timestamp 1666464484
transform 1 0 7820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_81
timestamp 1666464484
transform 1 0 8556 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_89
timestamp 1666464484
transform 1 0 9292 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_97
timestamp 1666464484
transform 1 0 10028 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_105
timestamp 1666464484
transform 1 0 10764 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_109
timestamp 1666464484
transform 1 0 11132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1666464484
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_113
timestamp 1666464484
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_121
timestamp 1666464484
transform 1 0 12236 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_129
timestamp 1666464484
transform 1 0 12972 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_137
timestamp 1666464484
transform 1 0 13708 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_145
timestamp 1666464484
transform 1 0 14444 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_153
timestamp 1666464484
transform 1 0 15180 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_161
timestamp 1666464484
transform 1 0 15916 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_165
timestamp 1666464484
transform 1 0 16284 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1666464484
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_169
timestamp 1666464484
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_177
timestamp 1666464484
transform 1 0 17388 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_185
timestamp 1666464484
transform 1 0 18124 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_193
timestamp 1666464484
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_201
timestamp 1666464484
transform 1 0 19596 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_209
timestamp 1666464484
transform 1 0 20332 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_217
timestamp 1666464484
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1666464484
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1666464484
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_225
timestamp 1666464484
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_233
timestamp 1666464484
transform 1 0 22540 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_241
timestamp 1666464484
transform 1 0 23276 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_249
timestamp 1666464484
transform 1 0 24012 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_257
timestamp 1666464484
transform 1 0 24748 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_265
timestamp 1666464484
transform 1 0 25484 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_273
timestamp 1666464484
transform 1 0 26220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_277
timestamp 1666464484
transform 1 0 26588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1666464484
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_281
timestamp 1666464484
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_289
timestamp 1666464484
transform 1 0 27692 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_297
timestamp 1666464484
transform 1 0 28428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_305
timestamp 1666464484
transform 1 0 29164 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_313
timestamp 1666464484
transform 1 0 29900 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_321
timestamp 1666464484
transform 1 0 30636 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_329
timestamp 1666464484
transform 1 0 31372 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_333
timestamp 1666464484
transform 1 0 31740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1666464484
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_337
timestamp 1666464484
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_345
timestamp 1666464484
transform 1 0 32844 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_353
timestamp 1666464484
transform 1 0 33580 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_361
timestamp 1666464484
transform 1 0 34316 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_369
timestamp 1666464484
transform 1 0 35052 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_377
timestamp 1666464484
transform 1 0 35788 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_385
timestamp 1666464484
transform 1 0 36524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_389
timestamp 1666464484
transform 1 0 36892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1666464484
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_393
timestamp 1666464484
transform 1 0 37260 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_401
timestamp 1666464484
transform 1 0 37996 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_409
timestamp 1666464484
transform 1 0 38732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_417
timestamp 1666464484
transform 1 0 39468 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_425
timestamp 1666464484
transform 1 0 40204 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_433
timestamp 1666464484
transform 1 0 40940 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_441
timestamp 1666464484
transform 1 0 41676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_445
timestamp 1666464484
transform 1 0 42044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1666464484
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_449
timestamp 1666464484
transform 1 0 42412 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_457
timestamp 1666464484
transform 1 0 43148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_465
timestamp 1666464484
transform 1 0 43884 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_473
timestamp 1666464484
transform 1 0 44620 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_481
timestamp 1666464484
transform 1 0 45356 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_489
timestamp 1666464484
transform 1 0 46092 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_497
timestamp 1666464484
transform 1 0 46828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_501
timestamp 1666464484
transform 1 0 47196 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1666464484
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_505
timestamp 1666464484
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_513
timestamp 1666464484
transform 1 0 48300 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_521
timestamp 1666464484
transform 1 0 49036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_529
timestamp 1666464484
transform 1 0 49772 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_537
timestamp 1666464484
transform 1 0 50508 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_545
timestamp 1666464484
transform 1 0 51244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_553
timestamp 1666464484
transform 1 0 51980 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_557
timestamp 1666464484
transform 1 0 52348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1666464484
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_561
timestamp 1666464484
transform 1 0 52716 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_569
timestamp 1666464484
transform 1 0 53452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_577
timestamp 1666464484
transform 1 0 54188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_585
timestamp 1666464484
transform 1 0 54924 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_593
timestamp 1666464484
transform 1 0 55660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_29_601
timestamp 1666464484
transform 1 0 56396 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_609
timestamp 1666464484
transform 1 0 57132 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_613
timestamp 1666464484
transform 1 0 57500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1666464484
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_29_617
timestamp 1666464484
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_3
timestamp 1666464484
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_11
timestamp 1666464484
transform 1 0 2116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_19
timestamp 1666464484
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1666464484
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_29
timestamp 1666464484
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_37
timestamp 1666464484
transform 1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_45
timestamp 1666464484
transform 1 0 5244 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_53
timestamp 1666464484
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_61
timestamp 1666464484
transform 1 0 6716 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_69
timestamp 1666464484
transform 1 0 7452 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_77
timestamp 1666464484
transform 1 0 8188 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_81
timestamp 1666464484
transform 1 0 8556 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1666464484
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_85
timestamp 1666464484
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_93
timestamp 1666464484
transform 1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_101
timestamp 1666464484
transform 1 0 10396 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_109
timestamp 1666464484
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_117
timestamp 1666464484
transform 1 0 11868 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_125
timestamp 1666464484
transform 1 0 12604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_133
timestamp 1666464484
transform 1 0 13340 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_137
timestamp 1666464484
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1666464484
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_141
timestamp 1666464484
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_149
timestamp 1666464484
transform 1 0 14812 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_157
timestamp 1666464484
transform 1 0 15548 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_165
timestamp 1666464484
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_173
timestamp 1666464484
transform 1 0 17020 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_181
timestamp 1666464484
transform 1 0 17756 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_189
timestamp 1666464484
transform 1 0 18492 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_193
timestamp 1666464484
transform 1 0 18860 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1666464484
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_197
timestamp 1666464484
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_205
timestamp 1666464484
transform 1 0 19964 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_213
timestamp 1666464484
transform 1 0 20700 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_221
timestamp 1666464484
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_229
timestamp 1666464484
transform 1 0 22172 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_237
timestamp 1666464484
transform 1 0 22908 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_245
timestamp 1666464484
transform 1 0 23644 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_249
timestamp 1666464484
transform 1 0 24012 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1666464484
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_253
timestamp 1666464484
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_261
timestamp 1666464484
transform 1 0 25116 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_269
timestamp 1666464484
transform 1 0 25852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_277
timestamp 1666464484
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_285
timestamp 1666464484
transform 1 0 27324 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_293
timestamp 1666464484
transform 1 0 28060 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_301
timestamp 1666464484
transform 1 0 28796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_305
timestamp 1666464484
transform 1 0 29164 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1666464484
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_309
timestamp 1666464484
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_317
timestamp 1666464484
transform 1 0 30268 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_325
timestamp 1666464484
transform 1 0 31004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_333
timestamp 1666464484
transform 1 0 31740 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_341
timestamp 1666464484
transform 1 0 32476 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_349
timestamp 1666464484
transform 1 0 33212 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_357
timestamp 1666464484
transform 1 0 33948 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_361
timestamp 1666464484
transform 1 0 34316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1666464484
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_365
timestamp 1666464484
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_373
timestamp 1666464484
transform 1 0 35420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_381
timestamp 1666464484
transform 1 0 36156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_389
timestamp 1666464484
transform 1 0 36892 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_397
timestamp 1666464484
transform 1 0 37628 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_405
timestamp 1666464484
transform 1 0 38364 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_413
timestamp 1666464484
transform 1 0 39100 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_417
timestamp 1666464484
transform 1 0 39468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1666464484
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_421
timestamp 1666464484
transform 1 0 39836 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_429
timestamp 1666464484
transform 1 0 40572 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_437
timestamp 1666464484
transform 1 0 41308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_445
timestamp 1666464484
transform 1 0 42044 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_453
timestamp 1666464484
transform 1 0 42780 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_461
timestamp 1666464484
transform 1 0 43516 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_469
timestamp 1666464484
transform 1 0 44252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_473
timestamp 1666464484
transform 1 0 44620 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1666464484
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_477
timestamp 1666464484
transform 1 0 44988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_485
timestamp 1666464484
transform 1 0 45724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_493
timestamp 1666464484
transform 1 0 46460 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_501
timestamp 1666464484
transform 1 0 47196 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_509
timestamp 1666464484
transform 1 0 47932 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_517
timestamp 1666464484
transform 1 0 48668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_525
timestamp 1666464484
transform 1 0 49404 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_529
timestamp 1666464484
transform 1 0 49772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1666464484
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_533
timestamp 1666464484
transform 1 0 50140 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_541
timestamp 1666464484
transform 1 0 50876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_549
timestamp 1666464484
transform 1 0 51612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_557
timestamp 1666464484
transform 1 0 52348 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_565
timestamp 1666464484
transform 1 0 53084 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_573
timestamp 1666464484
transform 1 0 53820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_581
timestamp 1666464484
transform 1 0 54556 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_585
timestamp 1666464484
transform 1 0 54924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1666464484
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_30_589
timestamp 1666464484
transform 1 0 55292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_597
timestamp 1666464484
transform 1 0 56028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_605
timestamp 1666464484
transform 1 0 56764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_30_613
timestamp 1666464484
transform 1 0 57500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_30_621
timestamp 1666464484
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_31_3
timestamp 1666464484
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_11
timestamp 1666464484
transform 1 0 2116 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_19
timestamp 1666464484
transform 1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_27
timestamp 1666464484
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_35
timestamp 1666464484
transform 1 0 4324 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_43
timestamp 1666464484
transform 1 0 5060 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_51
timestamp 1666464484
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1666464484
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_57
timestamp 1666464484
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_65
timestamp 1666464484
transform 1 0 7084 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_73
timestamp 1666464484
transform 1 0 7820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_81
timestamp 1666464484
transform 1 0 8556 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_89
timestamp 1666464484
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_97
timestamp 1666464484
transform 1 0 10028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_105
timestamp 1666464484
transform 1 0 10764 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1666464484
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1666464484
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_113
timestamp 1666464484
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_121
timestamp 1666464484
transform 1 0 12236 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_129
timestamp 1666464484
transform 1 0 12972 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_137
timestamp 1666464484
transform 1 0 13708 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_145
timestamp 1666464484
transform 1 0 14444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_153
timestamp 1666464484
transform 1 0 15180 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_161
timestamp 1666464484
transform 1 0 15916 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_165
timestamp 1666464484
transform 1 0 16284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1666464484
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_169
timestamp 1666464484
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_177
timestamp 1666464484
transform 1 0 17388 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_185
timestamp 1666464484
transform 1 0 18124 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_193
timestamp 1666464484
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_201
timestamp 1666464484
transform 1 0 19596 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_209
timestamp 1666464484
transform 1 0 20332 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_217
timestamp 1666464484
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1666464484
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1666464484
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_225
timestamp 1666464484
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_233
timestamp 1666464484
transform 1 0 22540 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_241
timestamp 1666464484
transform 1 0 23276 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_249
timestamp 1666464484
transform 1 0 24012 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_257
timestamp 1666464484
transform 1 0 24748 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_265
timestamp 1666464484
transform 1 0 25484 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_273
timestamp 1666464484
transform 1 0 26220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_277
timestamp 1666464484
transform 1 0 26588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1666464484
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_281
timestamp 1666464484
transform 1 0 26956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_289
timestamp 1666464484
transform 1 0 27692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_297
timestamp 1666464484
transform 1 0 28428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_305
timestamp 1666464484
transform 1 0 29164 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_313
timestamp 1666464484
transform 1 0 29900 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_321
timestamp 1666464484
transform 1 0 30636 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_329
timestamp 1666464484
transform 1 0 31372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_333
timestamp 1666464484
transform 1 0 31740 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1666464484
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_337
timestamp 1666464484
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_345
timestamp 1666464484
transform 1 0 32844 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_353
timestamp 1666464484
transform 1 0 33580 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_361
timestamp 1666464484
transform 1 0 34316 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_369
timestamp 1666464484
transform 1 0 35052 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_377
timestamp 1666464484
transform 1 0 35788 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_385
timestamp 1666464484
transform 1 0 36524 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_389
timestamp 1666464484
transform 1 0 36892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1666464484
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_393
timestamp 1666464484
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_401
timestamp 1666464484
transform 1 0 37996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_409
timestamp 1666464484
transform 1 0 38732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_417
timestamp 1666464484
transform 1 0 39468 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_425
timestamp 1666464484
transform 1 0 40204 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_433
timestamp 1666464484
transform 1 0 40940 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_441
timestamp 1666464484
transform 1 0 41676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_445
timestamp 1666464484
transform 1 0 42044 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1666464484
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_449
timestamp 1666464484
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_457
timestamp 1666464484
transform 1 0 43148 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_465
timestamp 1666464484
transform 1 0 43884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_473
timestamp 1666464484
transform 1 0 44620 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_481
timestamp 1666464484
transform 1 0 45356 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_489
timestamp 1666464484
transform 1 0 46092 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_497
timestamp 1666464484
transform 1 0 46828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_501
timestamp 1666464484
transform 1 0 47196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1666464484
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_505
timestamp 1666464484
transform 1 0 47564 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_513
timestamp 1666464484
transform 1 0 48300 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_521
timestamp 1666464484
transform 1 0 49036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_529
timestamp 1666464484
transform 1 0 49772 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_537
timestamp 1666464484
transform 1 0 50508 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_545
timestamp 1666464484
transform 1 0 51244 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_553
timestamp 1666464484
transform 1 0 51980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_557
timestamp 1666464484
transform 1 0 52348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1666464484
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_561
timestamp 1666464484
transform 1 0 52716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_569
timestamp 1666464484
transform 1 0 53452 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_577
timestamp 1666464484
transform 1 0 54188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_585
timestamp 1666464484
transform 1 0 54924 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_593
timestamp 1666464484
transform 1 0 55660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_31_601
timestamp 1666464484
transform 1 0 56396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_609
timestamp 1666464484
transform 1 0 57132 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_613
timestamp 1666464484
transform 1 0 57500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1666464484
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_617
timestamp 1666464484
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_3
timestamp 1666464484
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_11
timestamp 1666464484
transform 1 0 2116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_19
timestamp 1666464484
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1666464484
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_29
timestamp 1666464484
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_37
timestamp 1666464484
transform 1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_45
timestamp 1666464484
transform 1 0 5244 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_53
timestamp 1666464484
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_61
timestamp 1666464484
transform 1 0 6716 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_69
timestamp 1666464484
transform 1 0 7452 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_77
timestamp 1666464484
transform 1 0 8188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_81
timestamp 1666464484
transform 1 0 8556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1666464484
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_85
timestamp 1666464484
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_93
timestamp 1666464484
transform 1 0 9660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_101
timestamp 1666464484
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_109
timestamp 1666464484
transform 1 0 11132 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_117
timestamp 1666464484
transform 1 0 11868 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_125
timestamp 1666464484
transform 1 0 12604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_133
timestamp 1666464484
transform 1 0 13340 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_137
timestamp 1666464484
transform 1 0 13708 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1666464484
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_141
timestamp 1666464484
transform 1 0 14076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_149
timestamp 1666464484
transform 1 0 14812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_157
timestamp 1666464484
transform 1 0 15548 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_165
timestamp 1666464484
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_173
timestamp 1666464484
transform 1 0 17020 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_181
timestamp 1666464484
transform 1 0 17756 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_189
timestamp 1666464484
transform 1 0 18492 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_193
timestamp 1666464484
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1666464484
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_197
timestamp 1666464484
transform 1 0 19228 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_205
timestamp 1666464484
transform 1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_213
timestamp 1666464484
transform 1 0 20700 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_221
timestamp 1666464484
transform 1 0 21436 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_229
timestamp 1666464484
transform 1 0 22172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_237
timestamp 1666464484
transform 1 0 22908 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_245
timestamp 1666464484
transform 1 0 23644 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_249
timestamp 1666464484
transform 1 0 24012 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1666464484
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_253
timestamp 1666464484
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_261
timestamp 1666464484
transform 1 0 25116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_269
timestamp 1666464484
transform 1 0 25852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_277
timestamp 1666464484
transform 1 0 26588 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_285
timestamp 1666464484
transform 1 0 27324 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_293
timestamp 1666464484
transform 1 0 28060 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_301
timestamp 1666464484
transform 1 0 28796 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_305
timestamp 1666464484
transform 1 0 29164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1666464484
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_309
timestamp 1666464484
transform 1 0 29532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_317
timestamp 1666464484
transform 1 0 30268 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_325
timestamp 1666464484
transform 1 0 31004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_333
timestamp 1666464484
transform 1 0 31740 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_341
timestamp 1666464484
transform 1 0 32476 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_349
timestamp 1666464484
transform 1 0 33212 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_357
timestamp 1666464484
transform 1 0 33948 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_361
timestamp 1666464484
transform 1 0 34316 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1666464484
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_365
timestamp 1666464484
transform 1 0 34684 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_373
timestamp 1666464484
transform 1 0 35420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_381
timestamp 1666464484
transform 1 0 36156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_389
timestamp 1666464484
transform 1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_397
timestamp 1666464484
transform 1 0 37628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_405
timestamp 1666464484
transform 1 0 38364 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_413
timestamp 1666464484
transform 1 0 39100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_417
timestamp 1666464484
transform 1 0 39468 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1666464484
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_421
timestamp 1666464484
transform 1 0 39836 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_429
timestamp 1666464484
transform 1 0 40572 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_437
timestamp 1666464484
transform 1 0 41308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_445
timestamp 1666464484
transform 1 0 42044 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_453
timestamp 1666464484
transform 1 0 42780 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_461
timestamp 1666464484
transform 1 0 43516 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_469
timestamp 1666464484
transform 1 0 44252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_473
timestamp 1666464484
transform 1 0 44620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1666464484
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_477
timestamp 1666464484
transform 1 0 44988 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_485
timestamp 1666464484
transform 1 0 45724 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_493
timestamp 1666464484
transform 1 0 46460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_501
timestamp 1666464484
transform 1 0 47196 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_509
timestamp 1666464484
transform 1 0 47932 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_517
timestamp 1666464484
transform 1 0 48668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_525
timestamp 1666464484
transform 1 0 49404 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_529
timestamp 1666464484
transform 1 0 49772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1666464484
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_533
timestamp 1666464484
transform 1 0 50140 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_541
timestamp 1666464484
transform 1 0 50876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_549
timestamp 1666464484
transform 1 0 51612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_557
timestamp 1666464484
transform 1 0 52348 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_565
timestamp 1666464484
transform 1 0 53084 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_573
timestamp 1666464484
transform 1 0 53820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_581
timestamp 1666464484
transform 1 0 54556 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_585
timestamp 1666464484
transform 1 0 54924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1666464484
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_589
timestamp 1666464484
transform 1 0 55292 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_597
timestamp 1666464484
transform 1 0 56028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_605
timestamp 1666464484
transform 1 0 56764 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_613
timestamp 1666464484
transform 1 0 57500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_621
timestamp 1666464484
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_33_3
timestamp 1666464484
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_11
timestamp 1666464484
transform 1 0 2116 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_19
timestamp 1666464484
transform 1 0 2852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_27
timestamp 1666464484
transform 1 0 3588 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_35
timestamp 1666464484
transform 1 0 4324 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_43
timestamp 1666464484
transform 1 0 5060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_51
timestamp 1666464484
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1666464484
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_57
timestamp 1666464484
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_65
timestamp 1666464484
transform 1 0 7084 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_73
timestamp 1666464484
transform 1 0 7820 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_81
timestamp 1666464484
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_89
timestamp 1666464484
transform 1 0 9292 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_97
timestamp 1666464484
transform 1 0 10028 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_105
timestamp 1666464484
transform 1 0 10764 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_109
timestamp 1666464484
transform 1 0 11132 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1666464484
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_113
timestamp 1666464484
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_121
timestamp 1666464484
transform 1 0 12236 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_129
timestamp 1666464484
transform 1 0 12972 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_137
timestamp 1666464484
transform 1 0 13708 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_145
timestamp 1666464484
transform 1 0 14444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_153
timestamp 1666464484
transform 1 0 15180 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_161
timestamp 1666464484
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_165
timestamp 1666464484
transform 1 0 16284 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1666464484
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_169
timestamp 1666464484
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_177
timestamp 1666464484
transform 1 0 17388 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_185
timestamp 1666464484
transform 1 0 18124 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_193
timestamp 1666464484
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_201
timestamp 1666464484
transform 1 0 19596 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_209
timestamp 1666464484
transform 1 0 20332 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_217
timestamp 1666464484
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1666464484
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1666464484
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_225
timestamp 1666464484
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_233
timestamp 1666464484
transform 1 0 22540 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_241
timestamp 1666464484
transform 1 0 23276 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_249
timestamp 1666464484
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_257
timestamp 1666464484
transform 1 0 24748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_265
timestamp 1666464484
transform 1 0 25484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_273
timestamp 1666464484
transform 1 0 26220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_277
timestamp 1666464484
transform 1 0 26588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1666464484
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_281
timestamp 1666464484
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_289
timestamp 1666464484
transform 1 0 27692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_297
timestamp 1666464484
transform 1 0 28428 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_305
timestamp 1666464484
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_313
timestamp 1666464484
transform 1 0 29900 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_321
timestamp 1666464484
transform 1 0 30636 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_329
timestamp 1666464484
transform 1 0 31372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_333
timestamp 1666464484
transform 1 0 31740 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1666464484
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_337
timestamp 1666464484
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_345
timestamp 1666464484
transform 1 0 32844 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_353
timestamp 1666464484
transform 1 0 33580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_361
timestamp 1666464484
transform 1 0 34316 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_369
timestamp 1666464484
transform 1 0 35052 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_377
timestamp 1666464484
transform 1 0 35788 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_385
timestamp 1666464484
transform 1 0 36524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_389
timestamp 1666464484
transform 1 0 36892 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1666464484
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_393
timestamp 1666464484
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_401
timestamp 1666464484
transform 1 0 37996 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_409
timestamp 1666464484
transform 1 0 38732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_417
timestamp 1666464484
transform 1 0 39468 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_425
timestamp 1666464484
transform 1 0 40204 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_433
timestamp 1666464484
transform 1 0 40940 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_441
timestamp 1666464484
transform 1 0 41676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_445
timestamp 1666464484
transform 1 0 42044 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1666464484
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_449
timestamp 1666464484
transform 1 0 42412 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_457
timestamp 1666464484
transform 1 0 43148 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_465
timestamp 1666464484
transform 1 0 43884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_473
timestamp 1666464484
transform 1 0 44620 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_481
timestamp 1666464484
transform 1 0 45356 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_489
timestamp 1666464484
transform 1 0 46092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_497
timestamp 1666464484
transform 1 0 46828 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_501
timestamp 1666464484
transform 1 0 47196 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1666464484
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_505
timestamp 1666464484
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_513
timestamp 1666464484
transform 1 0 48300 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_521
timestamp 1666464484
transform 1 0 49036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_529
timestamp 1666464484
transform 1 0 49772 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_537
timestamp 1666464484
transform 1 0 50508 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_545
timestamp 1666464484
transform 1 0 51244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_553
timestamp 1666464484
transform 1 0 51980 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_557
timestamp 1666464484
transform 1 0 52348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1666464484
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_561
timestamp 1666464484
transform 1 0 52716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_569
timestamp 1666464484
transform 1 0 53452 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_577
timestamp 1666464484
transform 1 0 54188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_585
timestamp 1666464484
transform 1 0 54924 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_593
timestamp 1666464484
transform 1 0 55660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_33_601
timestamp 1666464484
transform 1 0 56396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_33_609
timestamp 1666464484
transform 1 0 57132 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_613
timestamp 1666464484
transform 1 0 57500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1666464484
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_33_617
timestamp 1666464484
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_3
timestamp 1666464484
transform 1 0 1380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_11
timestamp 1666464484
transform 1 0 2116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_19
timestamp 1666464484
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1666464484
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_29
timestamp 1666464484
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_37
timestamp 1666464484
transform 1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_45
timestamp 1666464484
transform 1 0 5244 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_53
timestamp 1666464484
transform 1 0 5980 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_61
timestamp 1666464484
transform 1 0 6716 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_69
timestamp 1666464484
transform 1 0 7452 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_77
timestamp 1666464484
transform 1 0 8188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_81
timestamp 1666464484
transform 1 0 8556 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1666464484
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_85
timestamp 1666464484
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_93
timestamp 1666464484
transform 1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_101
timestamp 1666464484
transform 1 0 10396 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_109
timestamp 1666464484
transform 1 0 11132 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_117
timestamp 1666464484
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_125
timestamp 1666464484
transform 1 0 12604 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_133
timestamp 1666464484
transform 1 0 13340 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_137
timestamp 1666464484
transform 1 0 13708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1666464484
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_141
timestamp 1666464484
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_149
timestamp 1666464484
transform 1 0 14812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_157
timestamp 1666464484
transform 1 0 15548 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_165
timestamp 1666464484
transform 1 0 16284 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_173
timestamp 1666464484
transform 1 0 17020 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_181
timestamp 1666464484
transform 1 0 17756 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_189
timestamp 1666464484
transform 1 0 18492 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_193
timestamp 1666464484
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1666464484
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_197
timestamp 1666464484
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_205
timestamp 1666464484
transform 1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_213
timestamp 1666464484
transform 1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_221
timestamp 1666464484
transform 1 0 21436 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_229
timestamp 1666464484
transform 1 0 22172 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_237
timestamp 1666464484
transform 1 0 22908 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_245
timestamp 1666464484
transform 1 0 23644 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_249
timestamp 1666464484
transform 1 0 24012 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1666464484
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_253
timestamp 1666464484
transform 1 0 24380 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_261
timestamp 1666464484
transform 1 0 25116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_269
timestamp 1666464484
transform 1 0 25852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_277
timestamp 1666464484
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_285
timestamp 1666464484
transform 1 0 27324 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_293
timestamp 1666464484
transform 1 0 28060 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_301
timestamp 1666464484
transform 1 0 28796 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_305
timestamp 1666464484
transform 1 0 29164 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1666464484
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_309
timestamp 1666464484
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_317
timestamp 1666464484
transform 1 0 30268 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_325
timestamp 1666464484
transform 1 0 31004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_333
timestamp 1666464484
transform 1 0 31740 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_341
timestamp 1666464484
transform 1 0 32476 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_349
timestamp 1666464484
transform 1 0 33212 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_357
timestamp 1666464484
transform 1 0 33948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_361
timestamp 1666464484
transform 1 0 34316 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1666464484
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_365
timestamp 1666464484
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_373
timestamp 1666464484
transform 1 0 35420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_381
timestamp 1666464484
transform 1 0 36156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_389
timestamp 1666464484
transform 1 0 36892 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_397
timestamp 1666464484
transform 1 0 37628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_405
timestamp 1666464484
transform 1 0 38364 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_413
timestamp 1666464484
transform 1 0 39100 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_417
timestamp 1666464484
transform 1 0 39468 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1666464484
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_421
timestamp 1666464484
transform 1 0 39836 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_429
timestamp 1666464484
transform 1 0 40572 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_437
timestamp 1666464484
transform 1 0 41308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_445
timestamp 1666464484
transform 1 0 42044 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_453
timestamp 1666464484
transform 1 0 42780 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_461
timestamp 1666464484
transform 1 0 43516 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_469
timestamp 1666464484
transform 1 0 44252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_473
timestamp 1666464484
transform 1 0 44620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1666464484
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_477
timestamp 1666464484
transform 1 0 44988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_485
timestamp 1666464484
transform 1 0 45724 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_493
timestamp 1666464484
transform 1 0 46460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_501
timestamp 1666464484
transform 1 0 47196 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_509
timestamp 1666464484
transform 1 0 47932 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_517
timestamp 1666464484
transform 1 0 48668 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_525
timestamp 1666464484
transform 1 0 49404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_529
timestamp 1666464484
transform 1 0 49772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1666464484
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_533
timestamp 1666464484
transform 1 0 50140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_541
timestamp 1666464484
transform 1 0 50876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_549
timestamp 1666464484
transform 1 0 51612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_557
timestamp 1666464484
transform 1 0 52348 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_565
timestamp 1666464484
transform 1 0 53084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_573
timestamp 1666464484
transform 1 0 53820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_581
timestamp 1666464484
transform 1 0 54556 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_585
timestamp 1666464484
transform 1 0 54924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1666464484
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_589
timestamp 1666464484
transform 1 0 55292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_597
timestamp 1666464484
transform 1 0 56028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_605
timestamp 1666464484
transform 1 0 56764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_34_613
timestamp 1666464484
transform 1 0 57500 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_34_621
timestamp 1666464484
transform 1 0 58236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_35_3
timestamp 1666464484
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_11
timestamp 1666464484
transform 1 0 2116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_19
timestamp 1666464484
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_27
timestamp 1666464484
transform 1 0 3588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_35
timestamp 1666464484
transform 1 0 4324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_43
timestamp 1666464484
transform 1 0 5060 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_51
timestamp 1666464484
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1666464484
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_57
timestamp 1666464484
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_65
timestamp 1666464484
transform 1 0 7084 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_73
timestamp 1666464484
transform 1 0 7820 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_81
timestamp 1666464484
transform 1 0 8556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_89
timestamp 1666464484
transform 1 0 9292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_97
timestamp 1666464484
transform 1 0 10028 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_105
timestamp 1666464484
transform 1 0 10764 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_109
timestamp 1666464484
transform 1 0 11132 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1666464484
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_113
timestamp 1666464484
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_121
timestamp 1666464484
transform 1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_129
timestamp 1666464484
transform 1 0 12972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_137
timestamp 1666464484
transform 1 0 13708 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_145
timestamp 1666464484
transform 1 0 14444 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_153
timestamp 1666464484
transform 1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_161
timestamp 1666464484
transform 1 0 15916 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_165
timestamp 1666464484
transform 1 0 16284 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1666464484
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_169
timestamp 1666464484
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_177
timestamp 1666464484
transform 1 0 17388 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_185
timestamp 1666464484
transform 1 0 18124 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_193
timestamp 1666464484
transform 1 0 18860 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_201
timestamp 1666464484
transform 1 0 19596 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_209
timestamp 1666464484
transform 1 0 20332 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_217
timestamp 1666464484
transform 1 0 21068 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_221
timestamp 1666464484
transform 1 0 21436 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1666464484
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_225
timestamp 1666464484
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_233
timestamp 1666464484
transform 1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_241
timestamp 1666464484
transform 1 0 23276 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_249
timestamp 1666464484
transform 1 0 24012 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_257
timestamp 1666464484
transform 1 0 24748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_265
timestamp 1666464484
transform 1 0 25484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_273
timestamp 1666464484
transform 1 0 26220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_277
timestamp 1666464484
transform 1 0 26588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1666464484
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_281
timestamp 1666464484
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_289
timestamp 1666464484
transform 1 0 27692 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_297
timestamp 1666464484
transform 1 0 28428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_305
timestamp 1666464484
transform 1 0 29164 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_313
timestamp 1666464484
transform 1 0 29900 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_321
timestamp 1666464484
transform 1 0 30636 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_329
timestamp 1666464484
transform 1 0 31372 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_333
timestamp 1666464484
transform 1 0 31740 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1666464484
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_337
timestamp 1666464484
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_345
timestamp 1666464484
transform 1 0 32844 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_353
timestamp 1666464484
transform 1 0 33580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_361
timestamp 1666464484
transform 1 0 34316 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_369
timestamp 1666464484
transform 1 0 35052 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_377
timestamp 1666464484
transform 1 0 35788 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_385
timestamp 1666464484
transform 1 0 36524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_389
timestamp 1666464484
transform 1 0 36892 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1666464484
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_393
timestamp 1666464484
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_401
timestamp 1666464484
transform 1 0 37996 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_409
timestamp 1666464484
transform 1 0 38732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_417
timestamp 1666464484
transform 1 0 39468 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_425
timestamp 1666464484
transform 1 0 40204 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_433
timestamp 1666464484
transform 1 0 40940 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_441
timestamp 1666464484
transform 1 0 41676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_445
timestamp 1666464484
transform 1 0 42044 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1666464484
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_449
timestamp 1666464484
transform 1 0 42412 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_457
timestamp 1666464484
transform 1 0 43148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_465
timestamp 1666464484
transform 1 0 43884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_473
timestamp 1666464484
transform 1 0 44620 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_481
timestamp 1666464484
transform 1 0 45356 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_489
timestamp 1666464484
transform 1 0 46092 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_497
timestamp 1666464484
transform 1 0 46828 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_501
timestamp 1666464484
transform 1 0 47196 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1666464484
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_505
timestamp 1666464484
transform 1 0 47564 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_513
timestamp 1666464484
transform 1 0 48300 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_521
timestamp 1666464484
transform 1 0 49036 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_529
timestamp 1666464484
transform 1 0 49772 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_537
timestamp 1666464484
transform 1 0 50508 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_545
timestamp 1666464484
transform 1 0 51244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_553
timestamp 1666464484
transform 1 0 51980 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_557
timestamp 1666464484
transform 1 0 52348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1666464484
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_561
timestamp 1666464484
transform 1 0 52716 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_569
timestamp 1666464484
transform 1 0 53452 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_577
timestamp 1666464484
transform 1 0 54188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_585
timestamp 1666464484
transform 1 0 54924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_593
timestamp 1666464484
transform 1 0 55660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_35_601
timestamp 1666464484
transform 1 0 56396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_609
timestamp 1666464484
transform 1 0 57132 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_613
timestamp 1666464484
transform 1 0 57500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1666464484
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_617
timestamp 1666464484
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_3
timestamp 1666464484
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_11
timestamp 1666464484
transform 1 0 2116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_19
timestamp 1666464484
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1666464484
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_29
timestamp 1666464484
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_37
timestamp 1666464484
transform 1 0 4508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_45
timestamp 1666464484
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_53
timestamp 1666464484
transform 1 0 5980 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_61
timestamp 1666464484
transform 1 0 6716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_69
timestamp 1666464484
transform 1 0 7452 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_77
timestamp 1666464484
transform 1 0 8188 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_81
timestamp 1666464484
transform 1 0 8556 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1666464484
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_85
timestamp 1666464484
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_93
timestamp 1666464484
transform 1 0 9660 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_101
timestamp 1666464484
transform 1 0 10396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_109
timestamp 1666464484
transform 1 0 11132 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_117
timestamp 1666464484
transform 1 0 11868 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_125
timestamp 1666464484
transform 1 0 12604 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_133
timestamp 1666464484
transform 1 0 13340 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_137
timestamp 1666464484
transform 1 0 13708 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1666464484
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_141
timestamp 1666464484
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_149
timestamp 1666464484
transform 1 0 14812 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_157
timestamp 1666464484
transform 1 0 15548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_165
timestamp 1666464484
transform 1 0 16284 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_173
timestamp 1666464484
transform 1 0 17020 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_181
timestamp 1666464484
transform 1 0 17756 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_189
timestamp 1666464484
transform 1 0 18492 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_193
timestamp 1666464484
transform 1 0 18860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1666464484
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_197
timestamp 1666464484
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_205
timestamp 1666464484
transform 1 0 19964 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_213
timestamp 1666464484
transform 1 0 20700 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_221
timestamp 1666464484
transform 1 0 21436 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_229
timestamp 1666464484
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_237
timestamp 1666464484
transform 1 0 22908 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_245
timestamp 1666464484
transform 1 0 23644 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_249
timestamp 1666464484
transform 1 0 24012 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1666464484
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_253
timestamp 1666464484
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_261
timestamp 1666464484
transform 1 0 25116 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_269
timestamp 1666464484
transform 1 0 25852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_277
timestamp 1666464484
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_285
timestamp 1666464484
transform 1 0 27324 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_293
timestamp 1666464484
transform 1 0 28060 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_301
timestamp 1666464484
transform 1 0 28796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_305
timestamp 1666464484
transform 1 0 29164 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1666464484
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_309
timestamp 1666464484
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_317
timestamp 1666464484
transform 1 0 30268 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_325
timestamp 1666464484
transform 1 0 31004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_333
timestamp 1666464484
transform 1 0 31740 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_341
timestamp 1666464484
transform 1 0 32476 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_349
timestamp 1666464484
transform 1 0 33212 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_357
timestamp 1666464484
transform 1 0 33948 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_361
timestamp 1666464484
transform 1 0 34316 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1666464484
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_365
timestamp 1666464484
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_373
timestamp 1666464484
transform 1 0 35420 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_381
timestamp 1666464484
transform 1 0 36156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_389
timestamp 1666464484
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_397
timestamp 1666464484
transform 1 0 37628 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_405
timestamp 1666464484
transform 1 0 38364 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_413
timestamp 1666464484
transform 1 0 39100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_417
timestamp 1666464484
transform 1 0 39468 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1666464484
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_421
timestamp 1666464484
transform 1 0 39836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_429
timestamp 1666464484
transform 1 0 40572 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_437
timestamp 1666464484
transform 1 0 41308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_445
timestamp 1666464484
transform 1 0 42044 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_453
timestamp 1666464484
transform 1 0 42780 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_461
timestamp 1666464484
transform 1 0 43516 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_469
timestamp 1666464484
transform 1 0 44252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_473
timestamp 1666464484
transform 1 0 44620 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1666464484
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_477
timestamp 1666464484
transform 1 0 44988 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_485
timestamp 1666464484
transform 1 0 45724 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_493
timestamp 1666464484
transform 1 0 46460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_501
timestamp 1666464484
transform 1 0 47196 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_509
timestamp 1666464484
transform 1 0 47932 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_517
timestamp 1666464484
transform 1 0 48668 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_525
timestamp 1666464484
transform 1 0 49404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_529
timestamp 1666464484
transform 1 0 49772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1666464484
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_533
timestamp 1666464484
transform 1 0 50140 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_541
timestamp 1666464484
transform 1 0 50876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_549
timestamp 1666464484
transform 1 0 51612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_557
timestamp 1666464484
transform 1 0 52348 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_565
timestamp 1666464484
transform 1 0 53084 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_573
timestamp 1666464484
transform 1 0 53820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_581
timestamp 1666464484
transform 1 0 54556 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_585
timestamp 1666464484
transform 1 0 54924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1666464484
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_589
timestamp 1666464484
transform 1 0 55292 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_597
timestamp 1666464484
transform 1 0 56028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_605
timestamp 1666464484
transform 1 0 56764 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_36_613
timestamp 1666464484
transform 1 0 57500 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_621
timestamp 1666464484
transform 1 0 58236 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_37_3
timestamp 1666464484
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_11
timestamp 1666464484
transform 1 0 2116 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_19
timestamp 1666464484
transform 1 0 2852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_27
timestamp 1666464484
transform 1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_35
timestamp 1666464484
transform 1 0 4324 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_43
timestamp 1666464484
transform 1 0 5060 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_51
timestamp 1666464484
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1666464484
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_57
timestamp 1666464484
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_65
timestamp 1666464484
transform 1 0 7084 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_73
timestamp 1666464484
transform 1 0 7820 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_81
timestamp 1666464484
transform 1 0 8556 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_89
timestamp 1666464484
transform 1 0 9292 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_97
timestamp 1666464484
transform 1 0 10028 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_105
timestamp 1666464484
transform 1 0 10764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_109
timestamp 1666464484
transform 1 0 11132 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1666464484
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_113
timestamp 1666464484
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_121
timestamp 1666464484
transform 1 0 12236 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_129
timestamp 1666464484
transform 1 0 12972 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_137
timestamp 1666464484
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_145
timestamp 1666464484
transform 1 0 14444 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_153
timestamp 1666464484
transform 1 0 15180 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_161
timestamp 1666464484
transform 1 0 15916 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_165
timestamp 1666464484
transform 1 0 16284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1666464484
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_169
timestamp 1666464484
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_177
timestamp 1666464484
transform 1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_185
timestamp 1666464484
transform 1 0 18124 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_193
timestamp 1666464484
transform 1 0 18860 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_201
timestamp 1666464484
transform 1 0 19596 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_209
timestamp 1666464484
transform 1 0 20332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_217
timestamp 1666464484
transform 1 0 21068 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_221
timestamp 1666464484
transform 1 0 21436 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1666464484
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_225
timestamp 1666464484
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_233
timestamp 1666464484
transform 1 0 22540 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_241
timestamp 1666464484
transform 1 0 23276 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_249
timestamp 1666464484
transform 1 0 24012 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_257
timestamp 1666464484
transform 1 0 24748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_265
timestamp 1666464484
transform 1 0 25484 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_273
timestamp 1666464484
transform 1 0 26220 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_277
timestamp 1666464484
transform 1 0 26588 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1666464484
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_281
timestamp 1666464484
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_289
timestamp 1666464484
transform 1 0 27692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_297
timestamp 1666464484
transform 1 0 28428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_305
timestamp 1666464484
transform 1 0 29164 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_313
timestamp 1666464484
transform 1 0 29900 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_321
timestamp 1666464484
transform 1 0 30636 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_329
timestamp 1666464484
transform 1 0 31372 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_333
timestamp 1666464484
transform 1 0 31740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1666464484
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_337
timestamp 1666464484
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_345
timestamp 1666464484
transform 1 0 32844 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_353
timestamp 1666464484
transform 1 0 33580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_361
timestamp 1666464484
transform 1 0 34316 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_369
timestamp 1666464484
transform 1 0 35052 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_377
timestamp 1666464484
transform 1 0 35788 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_385
timestamp 1666464484
transform 1 0 36524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_389
timestamp 1666464484
transform 1 0 36892 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1666464484
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_393
timestamp 1666464484
transform 1 0 37260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_401
timestamp 1666464484
transform 1 0 37996 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_409
timestamp 1666464484
transform 1 0 38732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_417
timestamp 1666464484
transform 1 0 39468 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_425
timestamp 1666464484
transform 1 0 40204 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_433
timestamp 1666464484
transform 1 0 40940 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_441
timestamp 1666464484
transform 1 0 41676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_445
timestamp 1666464484
transform 1 0 42044 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1666464484
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_449
timestamp 1666464484
transform 1 0 42412 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_457
timestamp 1666464484
transform 1 0 43148 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_465
timestamp 1666464484
transform 1 0 43884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_473
timestamp 1666464484
transform 1 0 44620 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_481
timestamp 1666464484
transform 1 0 45356 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_489
timestamp 1666464484
transform 1 0 46092 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_497
timestamp 1666464484
transform 1 0 46828 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_501
timestamp 1666464484
transform 1 0 47196 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1666464484
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_505
timestamp 1666464484
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_513
timestamp 1666464484
transform 1 0 48300 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_521
timestamp 1666464484
transform 1 0 49036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_529
timestamp 1666464484
transform 1 0 49772 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_537
timestamp 1666464484
transform 1 0 50508 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_545
timestamp 1666464484
transform 1 0 51244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_553
timestamp 1666464484
transform 1 0 51980 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_557
timestamp 1666464484
transform 1 0 52348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1666464484
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_561
timestamp 1666464484
transform 1 0 52716 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_569
timestamp 1666464484
transform 1 0 53452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_577
timestamp 1666464484
transform 1 0 54188 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_585
timestamp 1666464484
transform 1 0 54924 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_593
timestamp 1666464484
transform 1 0 55660 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_601
timestamp 1666464484
transform 1 0 56396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_609
timestamp 1666464484
transform 1 0 57132 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_613
timestamp 1666464484
transform 1 0 57500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1666464484
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_617
timestamp 1666464484
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_3
timestamp 1666464484
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_11
timestamp 1666464484
transform 1 0 2116 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_19
timestamp 1666464484
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1666464484
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_29
timestamp 1666464484
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_37
timestamp 1666464484
transform 1 0 4508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_45
timestamp 1666464484
transform 1 0 5244 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_53
timestamp 1666464484
transform 1 0 5980 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_61
timestamp 1666464484
transform 1 0 6716 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_69
timestamp 1666464484
transform 1 0 7452 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_77
timestamp 1666464484
transform 1 0 8188 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_81
timestamp 1666464484
transform 1 0 8556 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1666464484
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_85
timestamp 1666464484
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_93
timestamp 1666464484
transform 1 0 9660 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_101
timestamp 1666464484
transform 1 0 10396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_109
timestamp 1666464484
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_117
timestamp 1666464484
transform 1 0 11868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_125
timestamp 1666464484
transform 1 0 12604 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_133
timestamp 1666464484
transform 1 0 13340 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_137
timestamp 1666464484
transform 1 0 13708 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1666464484
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_141
timestamp 1666464484
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_149
timestamp 1666464484
transform 1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_157
timestamp 1666464484
transform 1 0 15548 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_165
timestamp 1666464484
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_173
timestamp 1666464484
transform 1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_181
timestamp 1666464484
transform 1 0 17756 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_189
timestamp 1666464484
transform 1 0 18492 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_193
timestamp 1666464484
transform 1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1666464484
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_197
timestamp 1666464484
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_205
timestamp 1666464484
transform 1 0 19964 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_213
timestamp 1666464484
transform 1 0 20700 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_221
timestamp 1666464484
transform 1 0 21436 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_229
timestamp 1666464484
transform 1 0 22172 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_237
timestamp 1666464484
transform 1 0 22908 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_245
timestamp 1666464484
transform 1 0 23644 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_249
timestamp 1666464484
transform 1 0 24012 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1666464484
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_253
timestamp 1666464484
transform 1 0 24380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_261
timestamp 1666464484
transform 1 0 25116 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_269
timestamp 1666464484
transform 1 0 25852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_277
timestamp 1666464484
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_285
timestamp 1666464484
transform 1 0 27324 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_293
timestamp 1666464484
transform 1 0 28060 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_301
timestamp 1666464484
transform 1 0 28796 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_305
timestamp 1666464484
transform 1 0 29164 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1666464484
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_309
timestamp 1666464484
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_317
timestamp 1666464484
transform 1 0 30268 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_325
timestamp 1666464484
transform 1 0 31004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_333
timestamp 1666464484
transform 1 0 31740 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_341
timestamp 1666464484
transform 1 0 32476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_349
timestamp 1666464484
transform 1 0 33212 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_357
timestamp 1666464484
transform 1 0 33948 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_361
timestamp 1666464484
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1666464484
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_365
timestamp 1666464484
transform 1 0 34684 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_373
timestamp 1666464484
transform 1 0 35420 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_381
timestamp 1666464484
transform 1 0 36156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_389
timestamp 1666464484
transform 1 0 36892 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_397
timestamp 1666464484
transform 1 0 37628 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_405
timestamp 1666464484
transform 1 0 38364 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_413
timestamp 1666464484
transform 1 0 39100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_417
timestamp 1666464484
transform 1 0 39468 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1666464484
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_421
timestamp 1666464484
transform 1 0 39836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_429
timestamp 1666464484
transform 1 0 40572 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_437
timestamp 1666464484
transform 1 0 41308 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_445
timestamp 1666464484
transform 1 0 42044 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_453
timestamp 1666464484
transform 1 0 42780 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_461
timestamp 1666464484
transform 1 0 43516 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_469
timestamp 1666464484
transform 1 0 44252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_473
timestamp 1666464484
transform 1 0 44620 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1666464484
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_477
timestamp 1666464484
transform 1 0 44988 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_485
timestamp 1666464484
transform 1 0 45724 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_493
timestamp 1666464484
transform 1 0 46460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_501
timestamp 1666464484
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_509
timestamp 1666464484
transform 1 0 47932 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_517
timestamp 1666464484
transform 1 0 48668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_525
timestamp 1666464484
transform 1 0 49404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_529
timestamp 1666464484
transform 1 0 49772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1666464484
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_533
timestamp 1666464484
transform 1 0 50140 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_541
timestamp 1666464484
transform 1 0 50876 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_549
timestamp 1666464484
transform 1 0 51612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_557
timestamp 1666464484
transform 1 0 52348 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_565
timestamp 1666464484
transform 1 0 53084 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_573
timestamp 1666464484
transform 1 0 53820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_581
timestamp 1666464484
transform 1 0 54556 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_585
timestamp 1666464484
transform 1 0 54924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1666464484
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_589
timestamp 1666464484
transform 1 0 55292 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_597
timestamp 1666464484
transform 1 0 56028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_605
timestamp 1666464484
transform 1 0 56764 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_613
timestamp 1666464484
transform 1 0 57500 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_38_621
timestamp 1666464484
transform 1 0 58236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_39_3
timestamp 1666464484
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_11
timestamp 1666464484
transform 1 0 2116 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_19
timestamp 1666464484
transform 1 0 2852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_27
timestamp 1666464484
transform 1 0 3588 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_35
timestamp 1666464484
transform 1 0 4324 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_43
timestamp 1666464484
transform 1 0 5060 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_51
timestamp 1666464484
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1666464484
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_57
timestamp 1666464484
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_65
timestamp 1666464484
transform 1 0 7084 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_73
timestamp 1666464484
transform 1 0 7820 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_81
timestamp 1666464484
transform 1 0 8556 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_89
timestamp 1666464484
transform 1 0 9292 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_97
timestamp 1666464484
transform 1 0 10028 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_105
timestamp 1666464484
transform 1 0 10764 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_109
timestamp 1666464484
transform 1 0 11132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1666464484
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_113
timestamp 1666464484
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_121
timestamp 1666464484
transform 1 0 12236 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_129
timestamp 1666464484
transform 1 0 12972 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_137
timestamp 1666464484
transform 1 0 13708 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_145
timestamp 1666464484
transform 1 0 14444 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_153
timestamp 1666464484
transform 1 0 15180 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_161
timestamp 1666464484
transform 1 0 15916 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_165
timestamp 1666464484
transform 1 0 16284 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1666464484
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_169
timestamp 1666464484
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_177
timestamp 1666464484
transform 1 0 17388 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_185
timestamp 1666464484
transform 1 0 18124 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_193
timestamp 1666464484
transform 1 0 18860 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_201
timestamp 1666464484
transform 1 0 19596 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_209
timestamp 1666464484
transform 1 0 20332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_217
timestamp 1666464484
transform 1 0 21068 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_221
timestamp 1666464484
transform 1 0 21436 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1666464484
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_225
timestamp 1666464484
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_233
timestamp 1666464484
transform 1 0 22540 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_241
timestamp 1666464484
transform 1 0 23276 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_249
timestamp 1666464484
transform 1 0 24012 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_257
timestamp 1666464484
transform 1 0 24748 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_265
timestamp 1666464484
transform 1 0 25484 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_273
timestamp 1666464484
transform 1 0 26220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_277
timestamp 1666464484
transform 1 0 26588 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1666464484
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_281
timestamp 1666464484
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_289
timestamp 1666464484
transform 1 0 27692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_297
timestamp 1666464484
transform 1 0 28428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_305
timestamp 1666464484
transform 1 0 29164 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_313
timestamp 1666464484
transform 1 0 29900 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_321
timestamp 1666464484
transform 1 0 30636 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_329
timestamp 1666464484
transform 1 0 31372 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_333
timestamp 1666464484
transform 1 0 31740 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1666464484
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_337
timestamp 1666464484
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_345
timestamp 1666464484
transform 1 0 32844 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_353
timestamp 1666464484
transform 1 0 33580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_361
timestamp 1666464484
transform 1 0 34316 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_369
timestamp 1666464484
transform 1 0 35052 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_377
timestamp 1666464484
transform 1 0 35788 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_385
timestamp 1666464484
transform 1 0 36524 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_389
timestamp 1666464484
transform 1 0 36892 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1666464484
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_393
timestamp 1666464484
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_401
timestamp 1666464484
transform 1 0 37996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_409
timestamp 1666464484
transform 1 0 38732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_417
timestamp 1666464484
transform 1 0 39468 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_425
timestamp 1666464484
transform 1 0 40204 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_433
timestamp 1666464484
transform 1 0 40940 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_441
timestamp 1666464484
transform 1 0 41676 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_445
timestamp 1666464484
transform 1 0 42044 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1666464484
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_449
timestamp 1666464484
transform 1 0 42412 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_457
timestamp 1666464484
transform 1 0 43148 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_465
timestamp 1666464484
transform 1 0 43884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_473
timestamp 1666464484
transform 1 0 44620 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_481
timestamp 1666464484
transform 1 0 45356 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_489
timestamp 1666464484
transform 1 0 46092 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_497
timestamp 1666464484
transform 1 0 46828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_501
timestamp 1666464484
transform 1 0 47196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1666464484
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_505
timestamp 1666464484
transform 1 0 47564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_513
timestamp 1666464484
transform 1 0 48300 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_521
timestamp 1666464484
transform 1 0 49036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_529
timestamp 1666464484
transform 1 0 49772 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_537
timestamp 1666464484
transform 1 0 50508 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_545
timestamp 1666464484
transform 1 0 51244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_553
timestamp 1666464484
transform 1 0 51980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_557
timestamp 1666464484
transform 1 0 52348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1666464484
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_561
timestamp 1666464484
transform 1 0 52716 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_569
timestamp 1666464484
transform 1 0 53452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_577
timestamp 1666464484
transform 1 0 54188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_585
timestamp 1666464484
transform 1 0 54924 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_593
timestamp 1666464484
transform 1 0 55660 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_39_601
timestamp 1666464484
transform 1 0 56396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_39_609
timestamp 1666464484
transform 1 0 57132 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_613
timestamp 1666464484
transform 1 0 57500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1666464484
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_617
timestamp 1666464484
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_3
timestamp 1666464484
transform 1 0 1380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_11
timestamp 1666464484
transform 1 0 2116 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_19
timestamp 1666464484
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1666464484
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_29
timestamp 1666464484
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_37
timestamp 1666464484
transform 1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_45
timestamp 1666464484
transform 1 0 5244 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_53
timestamp 1666464484
transform 1 0 5980 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_61
timestamp 1666464484
transform 1 0 6716 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_69
timestamp 1666464484
transform 1 0 7452 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_77
timestamp 1666464484
transform 1 0 8188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_81
timestamp 1666464484
transform 1 0 8556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1666464484
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_85
timestamp 1666464484
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_93
timestamp 1666464484
transform 1 0 9660 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_101
timestamp 1666464484
transform 1 0 10396 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_109
timestamp 1666464484
transform 1 0 11132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_117
timestamp 1666464484
transform 1 0 11868 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_125
timestamp 1666464484
transform 1 0 12604 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_133
timestamp 1666464484
transform 1 0 13340 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_137
timestamp 1666464484
transform 1 0 13708 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1666464484
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_141
timestamp 1666464484
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_149
timestamp 1666464484
transform 1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_157
timestamp 1666464484
transform 1 0 15548 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_165
timestamp 1666464484
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_173
timestamp 1666464484
transform 1 0 17020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_181
timestamp 1666464484
transform 1 0 17756 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_189
timestamp 1666464484
transform 1 0 18492 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_193
timestamp 1666464484
transform 1 0 18860 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1666464484
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_197
timestamp 1666464484
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_205
timestamp 1666464484
transform 1 0 19964 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_213
timestamp 1666464484
transform 1 0 20700 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_221
timestamp 1666464484
transform 1 0 21436 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_229
timestamp 1666464484
transform 1 0 22172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_237
timestamp 1666464484
transform 1 0 22908 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_245
timestamp 1666464484
transform 1 0 23644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_249
timestamp 1666464484
transform 1 0 24012 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1666464484
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_253
timestamp 1666464484
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_261
timestamp 1666464484
transform 1 0 25116 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_269
timestamp 1666464484
transform 1 0 25852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_277
timestamp 1666464484
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_285
timestamp 1666464484
transform 1 0 27324 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_293
timestamp 1666464484
transform 1 0 28060 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_301
timestamp 1666464484
transform 1 0 28796 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_305
timestamp 1666464484
transform 1 0 29164 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1666464484
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_309
timestamp 1666464484
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_317
timestamp 1666464484
transform 1 0 30268 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_325
timestamp 1666464484
transform 1 0 31004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_333
timestamp 1666464484
transform 1 0 31740 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_341
timestamp 1666464484
transform 1 0 32476 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_349
timestamp 1666464484
transform 1 0 33212 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_357
timestamp 1666464484
transform 1 0 33948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_361
timestamp 1666464484
transform 1 0 34316 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1666464484
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_365
timestamp 1666464484
transform 1 0 34684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_373
timestamp 1666464484
transform 1 0 35420 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_381
timestamp 1666464484
transform 1 0 36156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_389
timestamp 1666464484
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_397
timestamp 1666464484
transform 1 0 37628 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_405
timestamp 1666464484
transform 1 0 38364 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_413
timestamp 1666464484
transform 1 0 39100 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_417
timestamp 1666464484
transform 1 0 39468 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1666464484
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_421
timestamp 1666464484
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_429
timestamp 1666464484
transform 1 0 40572 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_437
timestamp 1666464484
transform 1 0 41308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_445
timestamp 1666464484
transform 1 0 42044 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_453
timestamp 1666464484
transform 1 0 42780 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_461
timestamp 1666464484
transform 1 0 43516 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_469
timestamp 1666464484
transform 1 0 44252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_473
timestamp 1666464484
transform 1 0 44620 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1666464484
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_477
timestamp 1666464484
transform 1 0 44988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_485
timestamp 1666464484
transform 1 0 45724 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_493
timestamp 1666464484
transform 1 0 46460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_501
timestamp 1666464484
transform 1 0 47196 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_509
timestamp 1666464484
transform 1 0 47932 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_517
timestamp 1666464484
transform 1 0 48668 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_525
timestamp 1666464484
transform 1 0 49404 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_529
timestamp 1666464484
transform 1 0 49772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1666464484
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_533
timestamp 1666464484
transform 1 0 50140 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_541
timestamp 1666464484
transform 1 0 50876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_549
timestamp 1666464484
transform 1 0 51612 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_557
timestamp 1666464484
transform 1 0 52348 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_565
timestamp 1666464484
transform 1 0 53084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_573
timestamp 1666464484
transform 1 0 53820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_581
timestamp 1666464484
transform 1 0 54556 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_585
timestamp 1666464484
transform 1 0 54924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1666464484
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_589
timestamp 1666464484
transform 1 0 55292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_597
timestamp 1666464484
transform 1 0 56028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_605
timestamp 1666464484
transform 1 0 56764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_40_613
timestamp 1666464484
transform 1 0 57500 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_621
timestamp 1666464484
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_41_3
timestamp 1666464484
transform 1 0 1380 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_11
timestamp 1666464484
transform 1 0 2116 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_19
timestamp 1666464484
transform 1 0 2852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_27
timestamp 1666464484
transform 1 0 3588 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_35
timestamp 1666464484
transform 1 0 4324 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_43
timestamp 1666464484
transform 1 0 5060 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_51
timestamp 1666464484
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1666464484
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_57
timestamp 1666464484
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_65
timestamp 1666464484
transform 1 0 7084 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_73
timestamp 1666464484
transform 1 0 7820 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_81
timestamp 1666464484
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_89
timestamp 1666464484
transform 1 0 9292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_97
timestamp 1666464484
transform 1 0 10028 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_105
timestamp 1666464484
transform 1 0 10764 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_109
timestamp 1666464484
transform 1 0 11132 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1666464484
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_113
timestamp 1666464484
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_121
timestamp 1666464484
transform 1 0 12236 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_129
timestamp 1666464484
transform 1 0 12972 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_137
timestamp 1666464484
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_145
timestamp 1666464484
transform 1 0 14444 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_153
timestamp 1666464484
transform 1 0 15180 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_161
timestamp 1666464484
transform 1 0 15916 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_165
timestamp 1666464484
transform 1 0 16284 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1666464484
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_169
timestamp 1666464484
transform 1 0 16652 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_177
timestamp 1666464484
transform 1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_185
timestamp 1666464484
transform 1 0 18124 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_193
timestamp 1666464484
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_201
timestamp 1666464484
transform 1 0 19596 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_209
timestamp 1666464484
transform 1 0 20332 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_217
timestamp 1666464484
transform 1 0 21068 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_221
timestamp 1666464484
transform 1 0 21436 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1666464484
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_225
timestamp 1666464484
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_233
timestamp 1666464484
transform 1 0 22540 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_241
timestamp 1666464484
transform 1 0 23276 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_249
timestamp 1666464484
transform 1 0 24012 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_257
timestamp 1666464484
transform 1 0 24748 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_265
timestamp 1666464484
transform 1 0 25484 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_273
timestamp 1666464484
transform 1 0 26220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_277
timestamp 1666464484
transform 1 0 26588 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1666464484
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_281
timestamp 1666464484
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_289
timestamp 1666464484
transform 1 0 27692 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_297
timestamp 1666464484
transform 1 0 28428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_305
timestamp 1666464484
transform 1 0 29164 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_313
timestamp 1666464484
transform 1 0 29900 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_321
timestamp 1666464484
transform 1 0 30636 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_329
timestamp 1666464484
transform 1 0 31372 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_333
timestamp 1666464484
transform 1 0 31740 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1666464484
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_337
timestamp 1666464484
transform 1 0 32108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_345
timestamp 1666464484
transform 1 0 32844 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_353
timestamp 1666464484
transform 1 0 33580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_361
timestamp 1666464484
transform 1 0 34316 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_369
timestamp 1666464484
transform 1 0 35052 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_377
timestamp 1666464484
transform 1 0 35788 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_385
timestamp 1666464484
transform 1 0 36524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_389
timestamp 1666464484
transform 1 0 36892 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1666464484
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_393
timestamp 1666464484
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_401
timestamp 1666464484
transform 1 0 37996 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_409
timestamp 1666464484
transform 1 0 38732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_417
timestamp 1666464484
transform 1 0 39468 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_425
timestamp 1666464484
transform 1 0 40204 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_433
timestamp 1666464484
transform 1 0 40940 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_441
timestamp 1666464484
transform 1 0 41676 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_445
timestamp 1666464484
transform 1 0 42044 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1666464484
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_449
timestamp 1666464484
transform 1 0 42412 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_457
timestamp 1666464484
transform 1 0 43148 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_465
timestamp 1666464484
transform 1 0 43884 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_473
timestamp 1666464484
transform 1 0 44620 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_481
timestamp 1666464484
transform 1 0 45356 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_489
timestamp 1666464484
transform 1 0 46092 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_497
timestamp 1666464484
transform 1 0 46828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_501
timestamp 1666464484
transform 1 0 47196 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1666464484
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_505
timestamp 1666464484
transform 1 0 47564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_513
timestamp 1666464484
transform 1 0 48300 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_521
timestamp 1666464484
transform 1 0 49036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_529
timestamp 1666464484
transform 1 0 49772 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_537
timestamp 1666464484
transform 1 0 50508 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_545
timestamp 1666464484
transform 1 0 51244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_553
timestamp 1666464484
transform 1 0 51980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_557
timestamp 1666464484
transform 1 0 52348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1666464484
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_561
timestamp 1666464484
transform 1 0 52716 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_569
timestamp 1666464484
transform 1 0 53452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_577
timestamp 1666464484
transform 1 0 54188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_585
timestamp 1666464484
transform 1 0 54924 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_593
timestamp 1666464484
transform 1 0 55660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_601
timestamp 1666464484
transform 1 0 56396 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_609
timestamp 1666464484
transform 1 0 57132 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_613
timestamp 1666464484
transform 1 0 57500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1666464484
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_617
timestamp 1666464484
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_3
timestamp 1666464484
transform 1 0 1380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_11
timestamp 1666464484
transform 1 0 2116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_19
timestamp 1666464484
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1666464484
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_29
timestamp 1666464484
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_37
timestamp 1666464484
transform 1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_45
timestamp 1666464484
transform 1 0 5244 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_53
timestamp 1666464484
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_61
timestamp 1666464484
transform 1 0 6716 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_69
timestamp 1666464484
transform 1 0 7452 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_77
timestamp 1666464484
transform 1 0 8188 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_81
timestamp 1666464484
transform 1 0 8556 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1666464484
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_85
timestamp 1666464484
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_93
timestamp 1666464484
transform 1 0 9660 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_101
timestamp 1666464484
transform 1 0 10396 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_109
timestamp 1666464484
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_117
timestamp 1666464484
transform 1 0 11868 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_125
timestamp 1666464484
transform 1 0 12604 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_133
timestamp 1666464484
transform 1 0 13340 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_137
timestamp 1666464484
transform 1 0 13708 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1666464484
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_141
timestamp 1666464484
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_149
timestamp 1666464484
transform 1 0 14812 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_157
timestamp 1666464484
transform 1 0 15548 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_165
timestamp 1666464484
transform 1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_173
timestamp 1666464484
transform 1 0 17020 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_181
timestamp 1666464484
transform 1 0 17756 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_189
timestamp 1666464484
transform 1 0 18492 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_193
timestamp 1666464484
transform 1 0 18860 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1666464484
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_197
timestamp 1666464484
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_205
timestamp 1666464484
transform 1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_213
timestamp 1666464484
transform 1 0 20700 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_221
timestamp 1666464484
transform 1 0 21436 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_229
timestamp 1666464484
transform 1 0 22172 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_237
timestamp 1666464484
transform 1 0 22908 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_245
timestamp 1666464484
transform 1 0 23644 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_249
timestamp 1666464484
transform 1 0 24012 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1666464484
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_253
timestamp 1666464484
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_261
timestamp 1666464484
transform 1 0 25116 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_269
timestamp 1666464484
transform 1 0 25852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_277
timestamp 1666464484
transform 1 0 26588 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_285
timestamp 1666464484
transform 1 0 27324 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_293
timestamp 1666464484
transform 1 0 28060 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_301
timestamp 1666464484
transform 1 0 28796 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_305
timestamp 1666464484
transform 1 0 29164 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1666464484
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_309
timestamp 1666464484
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_317
timestamp 1666464484
transform 1 0 30268 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_325
timestamp 1666464484
transform 1 0 31004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_333
timestamp 1666464484
transform 1 0 31740 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_341
timestamp 1666464484
transform 1 0 32476 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_349
timestamp 1666464484
transform 1 0 33212 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_357
timestamp 1666464484
transform 1 0 33948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_361
timestamp 1666464484
transform 1 0 34316 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1666464484
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_365
timestamp 1666464484
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_373
timestamp 1666464484
transform 1 0 35420 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_381
timestamp 1666464484
transform 1 0 36156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_389
timestamp 1666464484
transform 1 0 36892 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_397
timestamp 1666464484
transform 1 0 37628 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_405
timestamp 1666464484
transform 1 0 38364 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_413
timestamp 1666464484
transform 1 0 39100 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_417
timestamp 1666464484
transform 1 0 39468 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1666464484
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_421
timestamp 1666464484
transform 1 0 39836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_429
timestamp 1666464484
transform 1 0 40572 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_437
timestamp 1666464484
transform 1 0 41308 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_445
timestamp 1666464484
transform 1 0 42044 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_453
timestamp 1666464484
transform 1 0 42780 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_461
timestamp 1666464484
transform 1 0 43516 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_469
timestamp 1666464484
transform 1 0 44252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_473
timestamp 1666464484
transform 1 0 44620 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1666464484
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_477
timestamp 1666464484
transform 1 0 44988 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_485
timestamp 1666464484
transform 1 0 45724 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_493
timestamp 1666464484
transform 1 0 46460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_501
timestamp 1666464484
transform 1 0 47196 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_509
timestamp 1666464484
transform 1 0 47932 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_517
timestamp 1666464484
transform 1 0 48668 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_525
timestamp 1666464484
transform 1 0 49404 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_529
timestamp 1666464484
transform 1 0 49772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1666464484
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_533
timestamp 1666464484
transform 1 0 50140 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_541
timestamp 1666464484
transform 1 0 50876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_549
timestamp 1666464484
transform 1 0 51612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_557
timestamp 1666464484
transform 1 0 52348 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_565
timestamp 1666464484
transform 1 0 53084 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_573
timestamp 1666464484
transform 1 0 53820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_581
timestamp 1666464484
transform 1 0 54556 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_585
timestamp 1666464484
transform 1 0 54924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1666464484
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_42_589
timestamp 1666464484
transform 1 0 55292 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_597
timestamp 1666464484
transform 1 0 56028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_605
timestamp 1666464484
transform 1 0 56764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_42_613
timestamp 1666464484
transform 1 0 57500 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_42_621
timestamp 1666464484
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_43_3
timestamp 1666464484
transform 1 0 1380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_11
timestamp 1666464484
transform 1 0 2116 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_19
timestamp 1666464484
transform 1 0 2852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_27
timestamp 1666464484
transform 1 0 3588 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_35
timestamp 1666464484
transform 1 0 4324 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_43
timestamp 1666464484
transform 1 0 5060 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_51
timestamp 1666464484
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1666464484
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_57
timestamp 1666464484
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_65
timestamp 1666464484
transform 1 0 7084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_73
timestamp 1666464484
transform 1 0 7820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_81
timestamp 1666464484
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_89
timestamp 1666464484
transform 1 0 9292 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_97
timestamp 1666464484
transform 1 0 10028 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_105
timestamp 1666464484
transform 1 0 10764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_109
timestamp 1666464484
transform 1 0 11132 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1666464484
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_113
timestamp 1666464484
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_121
timestamp 1666464484
transform 1 0 12236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_129
timestamp 1666464484
transform 1 0 12972 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_137
timestamp 1666464484
transform 1 0 13708 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_145
timestamp 1666464484
transform 1 0 14444 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_153
timestamp 1666464484
transform 1 0 15180 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_161
timestamp 1666464484
transform 1 0 15916 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_165
timestamp 1666464484
transform 1 0 16284 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1666464484
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_169
timestamp 1666464484
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_177
timestamp 1666464484
transform 1 0 17388 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_185
timestamp 1666464484
transform 1 0 18124 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_193
timestamp 1666464484
transform 1 0 18860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_201
timestamp 1666464484
transform 1 0 19596 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_209
timestamp 1666464484
transform 1 0 20332 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_217
timestamp 1666464484
transform 1 0 21068 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_221
timestamp 1666464484
transform 1 0 21436 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1666464484
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_225
timestamp 1666464484
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_233
timestamp 1666464484
transform 1 0 22540 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_241
timestamp 1666464484
transform 1 0 23276 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_249
timestamp 1666464484
transform 1 0 24012 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_257
timestamp 1666464484
transform 1 0 24748 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_265
timestamp 1666464484
transform 1 0 25484 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_273
timestamp 1666464484
transform 1 0 26220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_277
timestamp 1666464484
transform 1 0 26588 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1666464484
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_281
timestamp 1666464484
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_289
timestamp 1666464484
transform 1 0 27692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_297
timestamp 1666464484
transform 1 0 28428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_305
timestamp 1666464484
transform 1 0 29164 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_313
timestamp 1666464484
transform 1 0 29900 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_321
timestamp 1666464484
transform 1 0 30636 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_329
timestamp 1666464484
transform 1 0 31372 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_333
timestamp 1666464484
transform 1 0 31740 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1666464484
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_337
timestamp 1666464484
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_345
timestamp 1666464484
transform 1 0 32844 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_353
timestamp 1666464484
transform 1 0 33580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_361
timestamp 1666464484
transform 1 0 34316 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_369
timestamp 1666464484
transform 1 0 35052 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_377
timestamp 1666464484
transform 1 0 35788 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_385
timestamp 1666464484
transform 1 0 36524 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_389
timestamp 1666464484
transform 1 0 36892 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1666464484
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_393
timestamp 1666464484
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_401
timestamp 1666464484
transform 1 0 37996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_409
timestamp 1666464484
transform 1 0 38732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_417
timestamp 1666464484
transform 1 0 39468 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_425
timestamp 1666464484
transform 1 0 40204 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_433
timestamp 1666464484
transform 1 0 40940 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_441
timestamp 1666464484
transform 1 0 41676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_445
timestamp 1666464484
transform 1 0 42044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1666464484
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_449
timestamp 1666464484
transform 1 0 42412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_457
timestamp 1666464484
transform 1 0 43148 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_465
timestamp 1666464484
transform 1 0 43884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_473
timestamp 1666464484
transform 1 0 44620 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_481
timestamp 1666464484
transform 1 0 45356 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_489
timestamp 1666464484
transform 1 0 46092 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_497
timestamp 1666464484
transform 1 0 46828 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_501
timestamp 1666464484
transform 1 0 47196 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1666464484
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_505
timestamp 1666464484
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_513
timestamp 1666464484
transform 1 0 48300 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_521
timestamp 1666464484
transform 1 0 49036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_529
timestamp 1666464484
transform 1 0 49772 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_537
timestamp 1666464484
transform 1 0 50508 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_545
timestamp 1666464484
transform 1 0 51244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_553
timestamp 1666464484
transform 1 0 51980 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_557
timestamp 1666464484
transform 1 0 52348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1666464484
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_561
timestamp 1666464484
transform 1 0 52716 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_569
timestamp 1666464484
transform 1 0 53452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_577
timestamp 1666464484
transform 1 0 54188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_585
timestamp 1666464484
transform 1 0 54924 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_593
timestamp 1666464484
transform 1 0 55660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_43_601
timestamp 1666464484
transform 1 0 56396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_609
timestamp 1666464484
transform 1 0 57132 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_613
timestamp 1666464484
transform 1 0 57500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1666464484
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_43_617
timestamp 1666464484
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_3
timestamp 1666464484
transform 1 0 1380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_11
timestamp 1666464484
transform 1 0 2116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_19
timestamp 1666464484
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1666464484
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_29
timestamp 1666464484
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_37
timestamp 1666464484
transform 1 0 4508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_45
timestamp 1666464484
transform 1 0 5244 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_53
timestamp 1666464484
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_61
timestamp 1666464484
transform 1 0 6716 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_69
timestamp 1666464484
transform 1 0 7452 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_77
timestamp 1666464484
transform 1 0 8188 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_81
timestamp 1666464484
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1666464484
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_85
timestamp 1666464484
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_93
timestamp 1666464484
transform 1 0 9660 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_101
timestamp 1666464484
transform 1 0 10396 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_109
timestamp 1666464484
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_117
timestamp 1666464484
transform 1 0 11868 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_125
timestamp 1666464484
transform 1 0 12604 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_133
timestamp 1666464484
transform 1 0 13340 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_137
timestamp 1666464484
transform 1 0 13708 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1666464484
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_141
timestamp 1666464484
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_149
timestamp 1666464484
transform 1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_157
timestamp 1666464484
transform 1 0 15548 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_165
timestamp 1666464484
transform 1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_173
timestamp 1666464484
transform 1 0 17020 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_181
timestamp 1666464484
transform 1 0 17756 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_189
timestamp 1666464484
transform 1 0 18492 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_193
timestamp 1666464484
transform 1 0 18860 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1666464484
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_197
timestamp 1666464484
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_205
timestamp 1666464484
transform 1 0 19964 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_213
timestamp 1666464484
transform 1 0 20700 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_221
timestamp 1666464484
transform 1 0 21436 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_229
timestamp 1666464484
transform 1 0 22172 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_237
timestamp 1666464484
transform 1 0 22908 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_245
timestamp 1666464484
transform 1 0 23644 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_249
timestamp 1666464484
transform 1 0 24012 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1666464484
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_253
timestamp 1666464484
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_261
timestamp 1666464484
transform 1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_269
timestamp 1666464484
transform 1 0 25852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_277
timestamp 1666464484
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_285
timestamp 1666464484
transform 1 0 27324 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_293
timestamp 1666464484
transform 1 0 28060 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_301
timestamp 1666464484
transform 1 0 28796 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_305
timestamp 1666464484
transform 1 0 29164 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1666464484
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_309
timestamp 1666464484
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_317
timestamp 1666464484
transform 1 0 30268 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_325
timestamp 1666464484
transform 1 0 31004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_333
timestamp 1666464484
transform 1 0 31740 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_341
timestamp 1666464484
transform 1 0 32476 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_349
timestamp 1666464484
transform 1 0 33212 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_357
timestamp 1666464484
transform 1 0 33948 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_361
timestamp 1666464484
transform 1 0 34316 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1666464484
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_365
timestamp 1666464484
transform 1 0 34684 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_373
timestamp 1666464484
transform 1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_381
timestamp 1666464484
transform 1 0 36156 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_389
timestamp 1666464484
transform 1 0 36892 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_397
timestamp 1666464484
transform 1 0 37628 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_405
timestamp 1666464484
transform 1 0 38364 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_413
timestamp 1666464484
transform 1 0 39100 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_417
timestamp 1666464484
transform 1 0 39468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1666464484
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_421
timestamp 1666464484
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_429
timestamp 1666464484
transform 1 0 40572 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_437
timestamp 1666464484
transform 1 0 41308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_445
timestamp 1666464484
transform 1 0 42044 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_453
timestamp 1666464484
transform 1 0 42780 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_461
timestamp 1666464484
transform 1 0 43516 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_469
timestamp 1666464484
transform 1 0 44252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_473
timestamp 1666464484
transform 1 0 44620 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1666464484
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_477
timestamp 1666464484
transform 1 0 44988 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_485
timestamp 1666464484
transform 1 0 45724 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_493
timestamp 1666464484
transform 1 0 46460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_501
timestamp 1666464484
transform 1 0 47196 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_509
timestamp 1666464484
transform 1 0 47932 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_517
timestamp 1666464484
transform 1 0 48668 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_525
timestamp 1666464484
transform 1 0 49404 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_529
timestamp 1666464484
transform 1 0 49772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1666464484
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_533
timestamp 1666464484
transform 1 0 50140 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_541
timestamp 1666464484
transform 1 0 50876 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_549
timestamp 1666464484
transform 1 0 51612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_557
timestamp 1666464484
transform 1 0 52348 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_565
timestamp 1666464484
transform 1 0 53084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_573
timestamp 1666464484
transform 1 0 53820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_581
timestamp 1666464484
transform 1 0 54556 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_585
timestamp 1666464484
transform 1 0 54924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1666464484
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_44_589
timestamp 1666464484
transform 1 0 55292 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_597
timestamp 1666464484
transform 1 0 56028 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_605
timestamp 1666464484
transform 1 0 56764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_44_613
timestamp 1666464484
transform 1 0 57500 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_621
timestamp 1666464484
transform 1 0 58236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_45_3
timestamp 1666464484
transform 1 0 1380 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_11
timestamp 1666464484
transform 1 0 2116 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_19
timestamp 1666464484
transform 1 0 2852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_27
timestamp 1666464484
transform 1 0 3588 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_35
timestamp 1666464484
transform 1 0 4324 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_43
timestamp 1666464484
transform 1 0 5060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_51
timestamp 1666464484
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1666464484
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_57
timestamp 1666464484
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_65
timestamp 1666464484
transform 1 0 7084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_73
timestamp 1666464484
transform 1 0 7820 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_81
timestamp 1666464484
transform 1 0 8556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_89
timestamp 1666464484
transform 1 0 9292 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_97
timestamp 1666464484
transform 1 0 10028 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_105
timestamp 1666464484
transform 1 0 10764 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_109
timestamp 1666464484
transform 1 0 11132 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1666464484
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_113
timestamp 1666464484
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_121
timestamp 1666464484
transform 1 0 12236 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_129
timestamp 1666464484
transform 1 0 12972 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_137
timestamp 1666464484
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_145
timestamp 1666464484
transform 1 0 14444 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_153
timestamp 1666464484
transform 1 0 15180 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_161
timestamp 1666464484
transform 1 0 15916 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_165
timestamp 1666464484
transform 1 0 16284 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1666464484
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_169
timestamp 1666464484
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_177
timestamp 1666464484
transform 1 0 17388 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_185
timestamp 1666464484
transform 1 0 18124 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_193
timestamp 1666464484
transform 1 0 18860 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_201
timestamp 1666464484
transform 1 0 19596 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_209
timestamp 1666464484
transform 1 0 20332 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_217
timestamp 1666464484
transform 1 0 21068 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_221
timestamp 1666464484
transform 1 0 21436 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1666464484
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_225
timestamp 1666464484
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_233
timestamp 1666464484
transform 1 0 22540 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_241
timestamp 1666464484
transform 1 0 23276 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_249
timestamp 1666464484
transform 1 0 24012 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_257
timestamp 1666464484
transform 1 0 24748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_265
timestamp 1666464484
transform 1 0 25484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_273
timestamp 1666464484
transform 1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_277
timestamp 1666464484
transform 1 0 26588 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1666464484
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_281
timestamp 1666464484
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_289
timestamp 1666464484
transform 1 0 27692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_297
timestamp 1666464484
transform 1 0 28428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_305
timestamp 1666464484
transform 1 0 29164 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_313
timestamp 1666464484
transform 1 0 29900 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_321
timestamp 1666464484
transform 1 0 30636 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_329
timestamp 1666464484
transform 1 0 31372 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_333
timestamp 1666464484
transform 1 0 31740 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1666464484
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_337
timestamp 1666464484
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_345
timestamp 1666464484
transform 1 0 32844 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_353
timestamp 1666464484
transform 1 0 33580 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_361
timestamp 1666464484
transform 1 0 34316 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_369
timestamp 1666464484
transform 1 0 35052 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_377
timestamp 1666464484
transform 1 0 35788 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_385
timestamp 1666464484
transform 1 0 36524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_389
timestamp 1666464484
transform 1 0 36892 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1666464484
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_393
timestamp 1666464484
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_401
timestamp 1666464484
transform 1 0 37996 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_409
timestamp 1666464484
transform 1 0 38732 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_417
timestamp 1666464484
transform 1 0 39468 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_425
timestamp 1666464484
transform 1 0 40204 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_433
timestamp 1666464484
transform 1 0 40940 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_441
timestamp 1666464484
transform 1 0 41676 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_445
timestamp 1666464484
transform 1 0 42044 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1666464484
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_449
timestamp 1666464484
transform 1 0 42412 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_457
timestamp 1666464484
transform 1 0 43148 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_465
timestamp 1666464484
transform 1 0 43884 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_473
timestamp 1666464484
transform 1 0 44620 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_481
timestamp 1666464484
transform 1 0 45356 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_489
timestamp 1666464484
transform 1 0 46092 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_497
timestamp 1666464484
transform 1 0 46828 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_501
timestamp 1666464484
transform 1 0 47196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1666464484
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_505
timestamp 1666464484
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_513
timestamp 1666464484
transform 1 0 48300 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_521
timestamp 1666464484
transform 1 0 49036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_529
timestamp 1666464484
transform 1 0 49772 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_537
timestamp 1666464484
transform 1 0 50508 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_545
timestamp 1666464484
transform 1 0 51244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_553
timestamp 1666464484
transform 1 0 51980 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_557
timestamp 1666464484
transform 1 0 52348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1666464484
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_561
timestamp 1666464484
transform 1 0 52716 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_569
timestamp 1666464484
transform 1 0 53452 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_577
timestamp 1666464484
transform 1 0 54188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_585
timestamp 1666464484
transform 1 0 54924 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_593
timestamp 1666464484
transform 1 0 55660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_45_601
timestamp 1666464484
transform 1 0 56396 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_609
timestamp 1666464484
transform 1 0 57132 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_613
timestamp 1666464484
transform 1 0 57500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1666464484
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_45_617
timestamp 1666464484
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_3
timestamp 1666464484
transform 1 0 1380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_11
timestamp 1666464484
transform 1 0 2116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_19
timestamp 1666464484
transform 1 0 2852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1666464484
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_29
timestamp 1666464484
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_37
timestamp 1666464484
transform 1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_45
timestamp 1666464484
transform 1 0 5244 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_53
timestamp 1666464484
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_61
timestamp 1666464484
transform 1 0 6716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_69
timestamp 1666464484
transform 1 0 7452 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_77
timestamp 1666464484
transform 1 0 8188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_81
timestamp 1666464484
transform 1 0 8556 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1666464484
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_85
timestamp 1666464484
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_93
timestamp 1666464484
transform 1 0 9660 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_101
timestamp 1666464484
transform 1 0 10396 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_109
timestamp 1666464484
transform 1 0 11132 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_117
timestamp 1666464484
transform 1 0 11868 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_125
timestamp 1666464484
transform 1 0 12604 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_133
timestamp 1666464484
transform 1 0 13340 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_137
timestamp 1666464484
transform 1 0 13708 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1666464484
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_141
timestamp 1666464484
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_149
timestamp 1666464484
transform 1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_157
timestamp 1666464484
transform 1 0 15548 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_165
timestamp 1666464484
transform 1 0 16284 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_173
timestamp 1666464484
transform 1 0 17020 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_181
timestamp 1666464484
transform 1 0 17756 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_189
timestamp 1666464484
transform 1 0 18492 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_193
timestamp 1666464484
transform 1 0 18860 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1666464484
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_197
timestamp 1666464484
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_205
timestamp 1666464484
transform 1 0 19964 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_213
timestamp 1666464484
transform 1 0 20700 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_221
timestamp 1666464484
transform 1 0 21436 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_229
timestamp 1666464484
transform 1 0 22172 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_237
timestamp 1666464484
transform 1 0 22908 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_245
timestamp 1666464484
transform 1 0 23644 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_249
timestamp 1666464484
transform 1 0 24012 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1666464484
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_253
timestamp 1666464484
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_261
timestamp 1666464484
transform 1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_269
timestamp 1666464484
transform 1 0 25852 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_277
timestamp 1666464484
transform 1 0 26588 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_285
timestamp 1666464484
transform 1 0 27324 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_293
timestamp 1666464484
transform 1 0 28060 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_301
timestamp 1666464484
transform 1 0 28796 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_305
timestamp 1666464484
transform 1 0 29164 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1666464484
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_309
timestamp 1666464484
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_317
timestamp 1666464484
transform 1 0 30268 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_325
timestamp 1666464484
transform 1 0 31004 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_333
timestamp 1666464484
transform 1 0 31740 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_341
timestamp 1666464484
transform 1 0 32476 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_349
timestamp 1666464484
transform 1 0 33212 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_357
timestamp 1666464484
transform 1 0 33948 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_361
timestamp 1666464484
transform 1 0 34316 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1666464484
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_365
timestamp 1666464484
transform 1 0 34684 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_373
timestamp 1666464484
transform 1 0 35420 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_381
timestamp 1666464484
transform 1 0 36156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_389
timestamp 1666464484
transform 1 0 36892 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_397
timestamp 1666464484
transform 1 0 37628 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_405
timestamp 1666464484
transform 1 0 38364 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_413
timestamp 1666464484
transform 1 0 39100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_417
timestamp 1666464484
transform 1 0 39468 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1666464484
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_421
timestamp 1666464484
transform 1 0 39836 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_429
timestamp 1666464484
transform 1 0 40572 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_437
timestamp 1666464484
transform 1 0 41308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_445
timestamp 1666464484
transform 1 0 42044 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_453
timestamp 1666464484
transform 1 0 42780 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_461
timestamp 1666464484
transform 1 0 43516 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_469
timestamp 1666464484
transform 1 0 44252 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_473
timestamp 1666464484
transform 1 0 44620 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1666464484
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_477
timestamp 1666464484
transform 1 0 44988 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_485
timestamp 1666464484
transform 1 0 45724 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_493
timestamp 1666464484
transform 1 0 46460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_501
timestamp 1666464484
transform 1 0 47196 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_509
timestamp 1666464484
transform 1 0 47932 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_517
timestamp 1666464484
transform 1 0 48668 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_525
timestamp 1666464484
transform 1 0 49404 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_529
timestamp 1666464484
transform 1 0 49772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1666464484
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_533
timestamp 1666464484
transform 1 0 50140 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_541
timestamp 1666464484
transform 1 0 50876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_549
timestamp 1666464484
transform 1 0 51612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_557
timestamp 1666464484
transform 1 0 52348 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_565
timestamp 1666464484
transform 1 0 53084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_573
timestamp 1666464484
transform 1 0 53820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_581
timestamp 1666464484
transform 1 0 54556 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_585
timestamp 1666464484
transform 1 0 54924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1666464484
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_46_589
timestamp 1666464484
transform 1 0 55292 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_597
timestamp 1666464484
transform 1 0 56028 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_605
timestamp 1666464484
transform 1 0 56764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_46_613
timestamp 1666464484
transform 1 0 57500 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_46_621
timestamp 1666464484
transform 1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_47_3
timestamp 1666464484
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_11
timestamp 1666464484
transform 1 0 2116 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_19
timestamp 1666464484
transform 1 0 2852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_27
timestamp 1666464484
transform 1 0 3588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_35
timestamp 1666464484
transform 1 0 4324 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_43
timestamp 1666464484
transform 1 0 5060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_51
timestamp 1666464484
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1666464484
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_57
timestamp 1666464484
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_65
timestamp 1666464484
transform 1 0 7084 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_73
timestamp 1666464484
transform 1 0 7820 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_81
timestamp 1666464484
transform 1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_89
timestamp 1666464484
transform 1 0 9292 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_97
timestamp 1666464484
transform 1 0 10028 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_105
timestamp 1666464484
transform 1 0 10764 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_109
timestamp 1666464484
transform 1 0 11132 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1666464484
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_113
timestamp 1666464484
transform 1 0 11500 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_121
timestamp 1666464484
transform 1 0 12236 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_129
timestamp 1666464484
transform 1 0 12972 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_137
timestamp 1666464484
transform 1 0 13708 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_145
timestamp 1666464484
transform 1 0 14444 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_153
timestamp 1666464484
transform 1 0 15180 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_161
timestamp 1666464484
transform 1 0 15916 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_165
timestamp 1666464484
transform 1 0 16284 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1666464484
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_169
timestamp 1666464484
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_177
timestamp 1666464484
transform 1 0 17388 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_185
timestamp 1666464484
transform 1 0 18124 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_193
timestamp 1666464484
transform 1 0 18860 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_201
timestamp 1666464484
transform 1 0 19596 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_209
timestamp 1666464484
transform 1 0 20332 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_217
timestamp 1666464484
transform 1 0 21068 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_221
timestamp 1666464484
transform 1 0 21436 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1666464484
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_225
timestamp 1666464484
transform 1 0 21804 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_233
timestamp 1666464484
transform 1 0 22540 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_241
timestamp 1666464484
transform 1 0 23276 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_249
timestamp 1666464484
transform 1 0 24012 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_257
timestamp 1666464484
transform 1 0 24748 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_265
timestamp 1666464484
transform 1 0 25484 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_273
timestamp 1666464484
transform 1 0 26220 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_277
timestamp 1666464484
transform 1 0 26588 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1666464484
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_281
timestamp 1666464484
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_289
timestamp 1666464484
transform 1 0 27692 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_297
timestamp 1666464484
transform 1 0 28428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_305
timestamp 1666464484
transform 1 0 29164 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_313
timestamp 1666464484
transform 1 0 29900 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_321
timestamp 1666464484
transform 1 0 30636 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_329
timestamp 1666464484
transform 1 0 31372 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_333
timestamp 1666464484
transform 1 0 31740 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1666464484
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_337
timestamp 1666464484
transform 1 0 32108 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_345
timestamp 1666464484
transform 1 0 32844 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_353
timestamp 1666464484
transform 1 0 33580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_361
timestamp 1666464484
transform 1 0 34316 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_369
timestamp 1666464484
transform 1 0 35052 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_377
timestamp 1666464484
transform 1 0 35788 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_385
timestamp 1666464484
transform 1 0 36524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_389
timestamp 1666464484
transform 1 0 36892 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1666464484
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_393
timestamp 1666464484
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_401
timestamp 1666464484
transform 1 0 37996 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_409
timestamp 1666464484
transform 1 0 38732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_417
timestamp 1666464484
transform 1 0 39468 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_425
timestamp 1666464484
transform 1 0 40204 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_433
timestamp 1666464484
transform 1 0 40940 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_441
timestamp 1666464484
transform 1 0 41676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_445
timestamp 1666464484
transform 1 0 42044 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1666464484
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_449
timestamp 1666464484
transform 1 0 42412 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_457
timestamp 1666464484
transform 1 0 43148 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_465
timestamp 1666464484
transform 1 0 43884 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_473
timestamp 1666464484
transform 1 0 44620 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_481
timestamp 1666464484
transform 1 0 45356 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_489
timestamp 1666464484
transform 1 0 46092 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_497
timestamp 1666464484
transform 1 0 46828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_501
timestamp 1666464484
transform 1 0 47196 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1666464484
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_505
timestamp 1666464484
transform 1 0 47564 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_513
timestamp 1666464484
transform 1 0 48300 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_521
timestamp 1666464484
transform 1 0 49036 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_529
timestamp 1666464484
transform 1 0 49772 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_537
timestamp 1666464484
transform 1 0 50508 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_545
timestamp 1666464484
transform 1 0 51244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_553
timestamp 1666464484
transform 1 0 51980 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_557
timestamp 1666464484
transform 1 0 52348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1666464484
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_561
timestamp 1666464484
transform 1 0 52716 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_569
timestamp 1666464484
transform 1 0 53452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_577
timestamp 1666464484
transform 1 0 54188 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_585
timestamp 1666464484
transform 1 0 54924 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_593
timestamp 1666464484
transform 1 0 55660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_601
timestamp 1666464484
transform 1 0 56396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_47_609
timestamp 1666464484
transform 1 0 57132 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_613
timestamp 1666464484
transform 1 0 57500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1666464484
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_617
timestamp 1666464484
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_3
timestamp 1666464484
transform 1 0 1380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_11
timestamp 1666464484
transform 1 0 2116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_19
timestamp 1666464484
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1666464484
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_29
timestamp 1666464484
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_37
timestamp 1666464484
transform 1 0 4508 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_45
timestamp 1666464484
transform 1 0 5244 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_53
timestamp 1666464484
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_61
timestamp 1666464484
transform 1 0 6716 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_69
timestamp 1666464484
transform 1 0 7452 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_77
timestamp 1666464484
transform 1 0 8188 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_81
timestamp 1666464484
transform 1 0 8556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1666464484
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_85
timestamp 1666464484
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_93
timestamp 1666464484
transform 1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_101
timestamp 1666464484
transform 1 0 10396 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_109
timestamp 1666464484
transform 1 0 11132 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_117
timestamp 1666464484
transform 1 0 11868 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_125
timestamp 1666464484
transform 1 0 12604 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_133
timestamp 1666464484
transform 1 0 13340 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_137
timestamp 1666464484
transform 1 0 13708 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1666464484
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_141
timestamp 1666464484
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_149
timestamp 1666464484
transform 1 0 14812 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_157
timestamp 1666464484
transform 1 0 15548 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_165
timestamp 1666464484
transform 1 0 16284 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_173
timestamp 1666464484
transform 1 0 17020 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_181
timestamp 1666464484
transform 1 0 17756 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_189
timestamp 1666464484
transform 1 0 18492 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_193
timestamp 1666464484
transform 1 0 18860 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1666464484
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_197
timestamp 1666464484
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_205
timestamp 1666464484
transform 1 0 19964 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_213
timestamp 1666464484
transform 1 0 20700 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_221
timestamp 1666464484
transform 1 0 21436 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_229
timestamp 1666464484
transform 1 0 22172 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_237
timestamp 1666464484
transform 1 0 22908 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_245
timestamp 1666464484
transform 1 0 23644 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_249
timestamp 1666464484
transform 1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1666464484
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_253
timestamp 1666464484
transform 1 0 24380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_261
timestamp 1666464484
transform 1 0 25116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_269
timestamp 1666464484
transform 1 0 25852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_277
timestamp 1666464484
transform 1 0 26588 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_285
timestamp 1666464484
transform 1 0 27324 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_293
timestamp 1666464484
transform 1 0 28060 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_301
timestamp 1666464484
transform 1 0 28796 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_305
timestamp 1666464484
transform 1 0 29164 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1666464484
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_309
timestamp 1666464484
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_317
timestamp 1666464484
transform 1 0 30268 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_325
timestamp 1666464484
transform 1 0 31004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_333
timestamp 1666464484
transform 1 0 31740 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_341
timestamp 1666464484
transform 1 0 32476 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_349
timestamp 1666464484
transform 1 0 33212 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_357
timestamp 1666464484
transform 1 0 33948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_361
timestamp 1666464484
transform 1 0 34316 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1666464484
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_365
timestamp 1666464484
transform 1 0 34684 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_373
timestamp 1666464484
transform 1 0 35420 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_381
timestamp 1666464484
transform 1 0 36156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_389
timestamp 1666464484
transform 1 0 36892 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_397
timestamp 1666464484
transform 1 0 37628 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_405
timestamp 1666464484
transform 1 0 38364 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_413
timestamp 1666464484
transform 1 0 39100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_417
timestamp 1666464484
transform 1 0 39468 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1666464484
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_421
timestamp 1666464484
transform 1 0 39836 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_429
timestamp 1666464484
transform 1 0 40572 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_437
timestamp 1666464484
transform 1 0 41308 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_445
timestamp 1666464484
transform 1 0 42044 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_453
timestamp 1666464484
transform 1 0 42780 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_461
timestamp 1666464484
transform 1 0 43516 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_469
timestamp 1666464484
transform 1 0 44252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_473
timestamp 1666464484
transform 1 0 44620 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1666464484
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_477
timestamp 1666464484
transform 1 0 44988 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_485
timestamp 1666464484
transform 1 0 45724 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_493
timestamp 1666464484
transform 1 0 46460 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_501
timestamp 1666464484
transform 1 0 47196 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_509
timestamp 1666464484
transform 1 0 47932 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_517
timestamp 1666464484
transform 1 0 48668 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_525
timestamp 1666464484
transform 1 0 49404 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_529
timestamp 1666464484
transform 1 0 49772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1666464484
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_533
timestamp 1666464484
transform 1 0 50140 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_541
timestamp 1666464484
transform 1 0 50876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_549
timestamp 1666464484
transform 1 0 51612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_557
timestamp 1666464484
transform 1 0 52348 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_565
timestamp 1666464484
transform 1 0 53084 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_573
timestamp 1666464484
transform 1 0 53820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_581
timestamp 1666464484
transform 1 0 54556 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_585
timestamp 1666464484
transform 1 0 54924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1666464484
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_48_589
timestamp 1666464484
transform 1 0 55292 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_597
timestamp 1666464484
transform 1 0 56028 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_605
timestamp 1666464484
transform 1 0 56764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_48_613
timestamp 1666464484
transform 1 0 57500 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_621
timestamp 1666464484
transform 1 0 58236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_49_3
timestamp 1666464484
transform 1 0 1380 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_11
timestamp 1666464484
transform 1 0 2116 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_19
timestamp 1666464484
transform 1 0 2852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_27
timestamp 1666464484
transform 1 0 3588 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_35
timestamp 1666464484
transform 1 0 4324 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_43
timestamp 1666464484
transform 1 0 5060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_51
timestamp 1666464484
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1666464484
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_57
timestamp 1666464484
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_65
timestamp 1666464484
transform 1 0 7084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_73
timestamp 1666464484
transform 1 0 7820 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_81
timestamp 1666464484
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_89
timestamp 1666464484
transform 1 0 9292 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_97
timestamp 1666464484
transform 1 0 10028 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_105
timestamp 1666464484
transform 1 0 10764 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_109
timestamp 1666464484
transform 1 0 11132 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1666464484
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_113
timestamp 1666464484
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_121
timestamp 1666464484
transform 1 0 12236 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_129
timestamp 1666464484
transform 1 0 12972 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_137
timestamp 1666464484
transform 1 0 13708 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_145
timestamp 1666464484
transform 1 0 14444 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_153
timestamp 1666464484
transform 1 0 15180 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_161
timestamp 1666464484
transform 1 0 15916 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_165
timestamp 1666464484
transform 1 0 16284 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1666464484
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_169
timestamp 1666464484
transform 1 0 16652 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_177
timestamp 1666464484
transform 1 0 17388 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_185
timestamp 1666464484
transform 1 0 18124 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_193
timestamp 1666464484
transform 1 0 18860 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_201
timestamp 1666464484
transform 1 0 19596 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_209
timestamp 1666464484
transform 1 0 20332 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_217
timestamp 1666464484
transform 1 0 21068 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_221
timestamp 1666464484
transform 1 0 21436 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1666464484
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_225
timestamp 1666464484
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_233
timestamp 1666464484
transform 1 0 22540 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_241
timestamp 1666464484
transform 1 0 23276 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_249
timestamp 1666464484
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_257
timestamp 1666464484
transform 1 0 24748 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_265
timestamp 1666464484
transform 1 0 25484 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_273
timestamp 1666464484
transform 1 0 26220 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_277
timestamp 1666464484
transform 1 0 26588 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1666464484
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_281
timestamp 1666464484
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_289
timestamp 1666464484
transform 1 0 27692 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_297
timestamp 1666464484
transform 1 0 28428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_305
timestamp 1666464484
transform 1 0 29164 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_313
timestamp 1666464484
transform 1 0 29900 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_321
timestamp 1666464484
transform 1 0 30636 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_329
timestamp 1666464484
transform 1 0 31372 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_333
timestamp 1666464484
transform 1 0 31740 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1666464484
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_337
timestamp 1666464484
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_345
timestamp 1666464484
transform 1 0 32844 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_353
timestamp 1666464484
transform 1 0 33580 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_361
timestamp 1666464484
transform 1 0 34316 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_369
timestamp 1666464484
transform 1 0 35052 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_377
timestamp 1666464484
transform 1 0 35788 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_385
timestamp 1666464484
transform 1 0 36524 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_389
timestamp 1666464484
transform 1 0 36892 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1666464484
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_393
timestamp 1666464484
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_401
timestamp 1666464484
transform 1 0 37996 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_409
timestamp 1666464484
transform 1 0 38732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_417
timestamp 1666464484
transform 1 0 39468 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_425
timestamp 1666464484
transform 1 0 40204 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_433
timestamp 1666464484
transform 1 0 40940 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_441
timestamp 1666464484
transform 1 0 41676 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_445
timestamp 1666464484
transform 1 0 42044 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1666464484
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_449
timestamp 1666464484
transform 1 0 42412 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_457
timestamp 1666464484
transform 1 0 43148 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_465
timestamp 1666464484
transform 1 0 43884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_473
timestamp 1666464484
transform 1 0 44620 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_481
timestamp 1666464484
transform 1 0 45356 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_489
timestamp 1666464484
transform 1 0 46092 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_497
timestamp 1666464484
transform 1 0 46828 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_501
timestamp 1666464484
transform 1 0 47196 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1666464484
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_505
timestamp 1666464484
transform 1 0 47564 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_513
timestamp 1666464484
transform 1 0 48300 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_521
timestamp 1666464484
transform 1 0 49036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_529
timestamp 1666464484
transform 1 0 49772 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_537
timestamp 1666464484
transform 1 0 50508 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_545
timestamp 1666464484
transform 1 0 51244 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_553
timestamp 1666464484
transform 1 0 51980 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_557
timestamp 1666464484
transform 1 0 52348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1666464484
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_561
timestamp 1666464484
transform 1 0 52716 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_569
timestamp 1666464484
transform 1 0 53452 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_577
timestamp 1666464484
transform 1 0 54188 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_585
timestamp 1666464484
transform 1 0 54924 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_593
timestamp 1666464484
transform 1 0 55660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_49_601
timestamp 1666464484
transform 1 0 56396 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_609
timestamp 1666464484
transform 1 0 57132 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_613
timestamp 1666464484
transform 1 0 57500 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1666464484
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_617
timestamp 1666464484
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_3
timestamp 1666464484
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_11
timestamp 1666464484
transform 1 0 2116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_19
timestamp 1666464484
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1666464484
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_29
timestamp 1666464484
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_37
timestamp 1666464484
transform 1 0 4508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_45
timestamp 1666464484
transform 1 0 5244 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_53
timestamp 1666464484
transform 1 0 5980 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_61
timestamp 1666464484
transform 1 0 6716 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_69
timestamp 1666464484
transform 1 0 7452 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_77
timestamp 1666464484
transform 1 0 8188 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_81
timestamp 1666464484
transform 1 0 8556 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1666464484
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_85
timestamp 1666464484
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_93
timestamp 1666464484
transform 1 0 9660 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_101
timestamp 1666464484
transform 1 0 10396 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_109
timestamp 1666464484
transform 1 0 11132 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_117
timestamp 1666464484
transform 1 0 11868 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_125
timestamp 1666464484
transform 1 0 12604 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_133
timestamp 1666464484
transform 1 0 13340 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_137
timestamp 1666464484
transform 1 0 13708 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1666464484
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_141
timestamp 1666464484
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_149
timestamp 1666464484
transform 1 0 14812 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_157
timestamp 1666464484
transform 1 0 15548 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_165
timestamp 1666464484
transform 1 0 16284 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_173
timestamp 1666464484
transform 1 0 17020 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_181
timestamp 1666464484
transform 1 0 17756 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_189
timestamp 1666464484
transform 1 0 18492 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_193
timestamp 1666464484
transform 1 0 18860 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1666464484
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_197
timestamp 1666464484
transform 1 0 19228 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_205
timestamp 1666464484
transform 1 0 19964 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_213
timestamp 1666464484
transform 1 0 20700 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_221
timestamp 1666464484
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_229
timestamp 1666464484
transform 1 0 22172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_237
timestamp 1666464484
transform 1 0 22908 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_245
timestamp 1666464484
transform 1 0 23644 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_249
timestamp 1666464484
transform 1 0 24012 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1666464484
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_253
timestamp 1666464484
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_261
timestamp 1666464484
transform 1 0 25116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_269
timestamp 1666464484
transform 1 0 25852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_277
timestamp 1666464484
transform 1 0 26588 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_285
timestamp 1666464484
transform 1 0 27324 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_293
timestamp 1666464484
transform 1 0 28060 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_301
timestamp 1666464484
transform 1 0 28796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_305
timestamp 1666464484
transform 1 0 29164 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1666464484
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_309
timestamp 1666464484
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_317
timestamp 1666464484
transform 1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_325
timestamp 1666464484
transform 1 0 31004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_333
timestamp 1666464484
transform 1 0 31740 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_341
timestamp 1666464484
transform 1 0 32476 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_349
timestamp 1666464484
transform 1 0 33212 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_357
timestamp 1666464484
transform 1 0 33948 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_361
timestamp 1666464484
transform 1 0 34316 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1666464484
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_365
timestamp 1666464484
transform 1 0 34684 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_373
timestamp 1666464484
transform 1 0 35420 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_381
timestamp 1666464484
transform 1 0 36156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_389
timestamp 1666464484
transform 1 0 36892 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_397
timestamp 1666464484
transform 1 0 37628 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_405
timestamp 1666464484
transform 1 0 38364 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_413
timestamp 1666464484
transform 1 0 39100 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_417
timestamp 1666464484
transform 1 0 39468 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1666464484
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_421
timestamp 1666464484
transform 1 0 39836 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_429
timestamp 1666464484
transform 1 0 40572 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_437
timestamp 1666464484
transform 1 0 41308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_445
timestamp 1666464484
transform 1 0 42044 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_453
timestamp 1666464484
transform 1 0 42780 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_461
timestamp 1666464484
transform 1 0 43516 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_469
timestamp 1666464484
transform 1 0 44252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_473
timestamp 1666464484
transform 1 0 44620 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1666464484
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_477
timestamp 1666464484
transform 1 0 44988 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_485
timestamp 1666464484
transform 1 0 45724 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_493
timestamp 1666464484
transform 1 0 46460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_501
timestamp 1666464484
transform 1 0 47196 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_509
timestamp 1666464484
transform 1 0 47932 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_517
timestamp 1666464484
transform 1 0 48668 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_525
timestamp 1666464484
transform 1 0 49404 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_529
timestamp 1666464484
transform 1 0 49772 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1666464484
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_533
timestamp 1666464484
transform 1 0 50140 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_541
timestamp 1666464484
transform 1 0 50876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_549
timestamp 1666464484
transform 1 0 51612 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_557
timestamp 1666464484
transform 1 0 52348 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_565
timestamp 1666464484
transform 1 0 53084 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_573
timestamp 1666464484
transform 1 0 53820 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_581
timestamp 1666464484
transform 1 0 54556 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_585
timestamp 1666464484
transform 1 0 54924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1666464484
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_50_589
timestamp 1666464484
transform 1 0 55292 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_597
timestamp 1666464484
transform 1 0 56028 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_605
timestamp 1666464484
transform 1 0 56764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_50_613
timestamp 1666464484
transform 1 0 57500 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_621
timestamp 1666464484
transform 1 0 58236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_51_3
timestamp 1666464484
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_11
timestamp 1666464484
transform 1 0 2116 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_19
timestamp 1666464484
transform 1 0 2852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_27
timestamp 1666464484
transform 1 0 3588 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_35
timestamp 1666464484
transform 1 0 4324 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_43
timestamp 1666464484
transform 1 0 5060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_51
timestamp 1666464484
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1666464484
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_57
timestamp 1666464484
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_65
timestamp 1666464484
transform 1 0 7084 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_73
timestamp 1666464484
transform 1 0 7820 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_81
timestamp 1666464484
transform 1 0 8556 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_89
timestamp 1666464484
transform 1 0 9292 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_97
timestamp 1666464484
transform 1 0 10028 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_105
timestamp 1666464484
transform 1 0 10764 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_109
timestamp 1666464484
transform 1 0 11132 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1666464484
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_113
timestamp 1666464484
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_121
timestamp 1666464484
transform 1 0 12236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_129
timestamp 1666464484
transform 1 0 12972 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_137
timestamp 1666464484
transform 1 0 13708 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_145
timestamp 1666464484
transform 1 0 14444 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_153
timestamp 1666464484
transform 1 0 15180 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_161
timestamp 1666464484
transform 1 0 15916 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_165
timestamp 1666464484
transform 1 0 16284 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1666464484
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_169
timestamp 1666464484
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_177
timestamp 1666464484
transform 1 0 17388 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_185
timestamp 1666464484
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_193
timestamp 1666464484
transform 1 0 18860 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_201
timestamp 1666464484
transform 1 0 19596 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_209
timestamp 1666464484
transform 1 0 20332 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_217
timestamp 1666464484
transform 1 0 21068 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_221
timestamp 1666464484
transform 1 0 21436 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1666464484
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_225
timestamp 1666464484
transform 1 0 21804 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_233
timestamp 1666464484
transform 1 0 22540 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_241
timestamp 1666464484
transform 1 0 23276 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_249
timestamp 1666464484
transform 1 0 24012 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_257
timestamp 1666464484
transform 1 0 24748 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_265
timestamp 1666464484
transform 1 0 25484 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_273
timestamp 1666464484
transform 1 0 26220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_277
timestamp 1666464484
transform 1 0 26588 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1666464484
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_281
timestamp 1666464484
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_289
timestamp 1666464484
transform 1 0 27692 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_297
timestamp 1666464484
transform 1 0 28428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_305
timestamp 1666464484
transform 1 0 29164 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_313
timestamp 1666464484
transform 1 0 29900 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_321
timestamp 1666464484
transform 1 0 30636 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_329
timestamp 1666464484
transform 1 0 31372 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_333
timestamp 1666464484
transform 1 0 31740 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1666464484
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_337
timestamp 1666464484
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_345
timestamp 1666464484
transform 1 0 32844 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_353
timestamp 1666464484
transform 1 0 33580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_361
timestamp 1666464484
transform 1 0 34316 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_369
timestamp 1666464484
transform 1 0 35052 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_377
timestamp 1666464484
transform 1 0 35788 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_385
timestamp 1666464484
transform 1 0 36524 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_389
timestamp 1666464484
transform 1 0 36892 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1666464484
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_393
timestamp 1666464484
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_401
timestamp 1666464484
transform 1 0 37996 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_409
timestamp 1666464484
transform 1 0 38732 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_417
timestamp 1666464484
transform 1 0 39468 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_425
timestamp 1666464484
transform 1 0 40204 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_433
timestamp 1666464484
transform 1 0 40940 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_441
timestamp 1666464484
transform 1 0 41676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_445
timestamp 1666464484
transform 1 0 42044 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1666464484
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_449
timestamp 1666464484
transform 1 0 42412 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_457
timestamp 1666464484
transform 1 0 43148 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_465
timestamp 1666464484
transform 1 0 43884 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_473
timestamp 1666464484
transform 1 0 44620 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_481
timestamp 1666464484
transform 1 0 45356 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_489
timestamp 1666464484
transform 1 0 46092 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_497
timestamp 1666464484
transform 1 0 46828 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_501
timestamp 1666464484
transform 1 0 47196 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1666464484
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_505
timestamp 1666464484
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_513
timestamp 1666464484
transform 1 0 48300 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_521
timestamp 1666464484
transform 1 0 49036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_529
timestamp 1666464484
transform 1 0 49772 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_537
timestamp 1666464484
transform 1 0 50508 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_545
timestamp 1666464484
transform 1 0 51244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_553
timestamp 1666464484
transform 1 0 51980 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_557
timestamp 1666464484
transform 1 0 52348 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1666464484
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_561
timestamp 1666464484
transform 1 0 52716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_569
timestamp 1666464484
transform 1 0 53452 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_577
timestamp 1666464484
transform 1 0 54188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_585
timestamp 1666464484
transform 1 0 54924 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_593
timestamp 1666464484
transform 1 0 55660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_51_601
timestamp 1666464484
transform 1 0 56396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_51_609
timestamp 1666464484
transform 1 0 57132 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_613
timestamp 1666464484
transform 1 0 57500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1666464484
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_617
timestamp 1666464484
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_3
timestamp 1666464484
transform 1 0 1380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_11
timestamp 1666464484
transform 1 0 2116 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_19
timestamp 1666464484
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1666464484
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_29
timestamp 1666464484
transform 1 0 3772 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_37
timestamp 1666464484
transform 1 0 4508 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_45
timestamp 1666464484
transform 1 0 5244 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_53
timestamp 1666464484
transform 1 0 5980 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_61
timestamp 1666464484
transform 1 0 6716 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_69
timestamp 1666464484
transform 1 0 7452 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_77
timestamp 1666464484
transform 1 0 8188 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_81
timestamp 1666464484
transform 1 0 8556 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1666464484
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_85
timestamp 1666464484
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_93
timestamp 1666464484
transform 1 0 9660 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_101
timestamp 1666464484
transform 1 0 10396 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_109
timestamp 1666464484
transform 1 0 11132 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_117
timestamp 1666464484
transform 1 0 11868 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_125
timestamp 1666464484
transform 1 0 12604 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_133
timestamp 1666464484
transform 1 0 13340 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_137
timestamp 1666464484
transform 1 0 13708 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1666464484
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_141
timestamp 1666464484
transform 1 0 14076 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_149
timestamp 1666464484
transform 1 0 14812 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_157
timestamp 1666464484
transform 1 0 15548 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_165
timestamp 1666464484
transform 1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_173
timestamp 1666464484
transform 1 0 17020 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_181
timestamp 1666464484
transform 1 0 17756 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_189
timestamp 1666464484
transform 1 0 18492 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_193
timestamp 1666464484
transform 1 0 18860 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1666464484
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_197
timestamp 1666464484
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_205
timestamp 1666464484
transform 1 0 19964 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_213
timestamp 1666464484
transform 1 0 20700 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_221
timestamp 1666464484
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_229
timestamp 1666464484
transform 1 0 22172 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_237
timestamp 1666464484
transform 1 0 22908 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_245
timestamp 1666464484
transform 1 0 23644 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_249
timestamp 1666464484
transform 1 0 24012 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1666464484
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_253
timestamp 1666464484
transform 1 0 24380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_261
timestamp 1666464484
transform 1 0 25116 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_269
timestamp 1666464484
transform 1 0 25852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_277
timestamp 1666464484
transform 1 0 26588 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_285
timestamp 1666464484
transform 1 0 27324 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_293
timestamp 1666464484
transform 1 0 28060 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_301
timestamp 1666464484
transform 1 0 28796 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_305
timestamp 1666464484
transform 1 0 29164 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1666464484
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_309
timestamp 1666464484
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_317
timestamp 1666464484
transform 1 0 30268 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_325
timestamp 1666464484
transform 1 0 31004 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_333
timestamp 1666464484
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_341
timestamp 1666464484
transform 1 0 32476 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_349
timestamp 1666464484
transform 1 0 33212 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_357
timestamp 1666464484
transform 1 0 33948 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_361
timestamp 1666464484
transform 1 0 34316 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1666464484
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_365
timestamp 1666464484
transform 1 0 34684 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_373
timestamp 1666464484
transform 1 0 35420 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_381
timestamp 1666464484
transform 1 0 36156 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_389
timestamp 1666464484
transform 1 0 36892 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_397
timestamp 1666464484
transform 1 0 37628 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_405
timestamp 1666464484
transform 1 0 38364 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_413
timestamp 1666464484
transform 1 0 39100 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_417
timestamp 1666464484
transform 1 0 39468 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1666464484
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_421
timestamp 1666464484
transform 1 0 39836 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_429
timestamp 1666464484
transform 1 0 40572 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_437
timestamp 1666464484
transform 1 0 41308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_445
timestamp 1666464484
transform 1 0 42044 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_453
timestamp 1666464484
transform 1 0 42780 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_461
timestamp 1666464484
transform 1 0 43516 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_469
timestamp 1666464484
transform 1 0 44252 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_473
timestamp 1666464484
transform 1 0 44620 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1666464484
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_477
timestamp 1666464484
transform 1 0 44988 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_485
timestamp 1666464484
transform 1 0 45724 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_493
timestamp 1666464484
transform 1 0 46460 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_501
timestamp 1666464484
transform 1 0 47196 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_509
timestamp 1666464484
transform 1 0 47932 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_517
timestamp 1666464484
transform 1 0 48668 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_525
timestamp 1666464484
transform 1 0 49404 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_529
timestamp 1666464484
transform 1 0 49772 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1666464484
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_533
timestamp 1666464484
transform 1 0 50140 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_541
timestamp 1666464484
transform 1 0 50876 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_549
timestamp 1666464484
transform 1 0 51612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_557
timestamp 1666464484
transform 1 0 52348 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_565
timestamp 1666464484
transform 1 0 53084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_573
timestamp 1666464484
transform 1 0 53820 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_581
timestamp 1666464484
transform 1 0 54556 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_585
timestamp 1666464484
transform 1 0 54924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1666464484
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_589
timestamp 1666464484
transform 1 0 55292 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_597
timestamp 1666464484
transform 1 0 56028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_605
timestamp 1666464484
transform 1 0 56764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_52_613
timestamp 1666464484
transform 1 0 57500 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_52_621
timestamp 1666464484
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_53_3
timestamp 1666464484
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_11
timestamp 1666464484
transform 1 0 2116 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_19
timestamp 1666464484
transform 1 0 2852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_27
timestamp 1666464484
transform 1 0 3588 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_35
timestamp 1666464484
transform 1 0 4324 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_43
timestamp 1666464484
transform 1 0 5060 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_51
timestamp 1666464484
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1666464484
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_57
timestamp 1666464484
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_65
timestamp 1666464484
transform 1 0 7084 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_73
timestamp 1666464484
transform 1 0 7820 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_81
timestamp 1666464484
transform 1 0 8556 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_89
timestamp 1666464484
transform 1 0 9292 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_97
timestamp 1666464484
transform 1 0 10028 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_105
timestamp 1666464484
transform 1 0 10764 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_109
timestamp 1666464484
transform 1 0 11132 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1666464484
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_113
timestamp 1666464484
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_121
timestamp 1666464484
transform 1 0 12236 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_129
timestamp 1666464484
transform 1 0 12972 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_137
timestamp 1666464484
transform 1 0 13708 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_145
timestamp 1666464484
transform 1 0 14444 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_153
timestamp 1666464484
transform 1 0 15180 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_161
timestamp 1666464484
transform 1 0 15916 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_165
timestamp 1666464484
transform 1 0 16284 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1666464484
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_169
timestamp 1666464484
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_177
timestamp 1666464484
transform 1 0 17388 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_185
timestamp 1666464484
transform 1 0 18124 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_193
timestamp 1666464484
transform 1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_201
timestamp 1666464484
transform 1 0 19596 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_209
timestamp 1666464484
transform 1 0 20332 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_217
timestamp 1666464484
transform 1 0 21068 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_221
timestamp 1666464484
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1666464484
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_225
timestamp 1666464484
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_233
timestamp 1666464484
transform 1 0 22540 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_241
timestamp 1666464484
transform 1 0 23276 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_249
timestamp 1666464484
transform 1 0 24012 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_257
timestamp 1666464484
transform 1 0 24748 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_265
timestamp 1666464484
transform 1 0 25484 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_273
timestamp 1666464484
transform 1 0 26220 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_277
timestamp 1666464484
transform 1 0 26588 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1666464484
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_281
timestamp 1666464484
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_289
timestamp 1666464484
transform 1 0 27692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_297
timestamp 1666464484
transform 1 0 28428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_305
timestamp 1666464484
transform 1 0 29164 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_313
timestamp 1666464484
transform 1 0 29900 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_321
timestamp 1666464484
transform 1 0 30636 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_329
timestamp 1666464484
transform 1 0 31372 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_333
timestamp 1666464484
transform 1 0 31740 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1666464484
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_337
timestamp 1666464484
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_345
timestamp 1666464484
transform 1 0 32844 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_353
timestamp 1666464484
transform 1 0 33580 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_361
timestamp 1666464484
transform 1 0 34316 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_369
timestamp 1666464484
transform 1 0 35052 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_377
timestamp 1666464484
transform 1 0 35788 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_385
timestamp 1666464484
transform 1 0 36524 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_389
timestamp 1666464484
transform 1 0 36892 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1666464484
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_393
timestamp 1666464484
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_401
timestamp 1666464484
transform 1 0 37996 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_409
timestamp 1666464484
transform 1 0 38732 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_417
timestamp 1666464484
transform 1 0 39468 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_425
timestamp 1666464484
transform 1 0 40204 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_433
timestamp 1666464484
transform 1 0 40940 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_441
timestamp 1666464484
transform 1 0 41676 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_445
timestamp 1666464484
transform 1 0 42044 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1666464484
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_449
timestamp 1666464484
transform 1 0 42412 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_457
timestamp 1666464484
transform 1 0 43148 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_465
timestamp 1666464484
transform 1 0 43884 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_473
timestamp 1666464484
transform 1 0 44620 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_481
timestamp 1666464484
transform 1 0 45356 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_489
timestamp 1666464484
transform 1 0 46092 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_497
timestamp 1666464484
transform 1 0 46828 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_501
timestamp 1666464484
transform 1 0 47196 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1666464484
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_505
timestamp 1666464484
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_513
timestamp 1666464484
transform 1 0 48300 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_521
timestamp 1666464484
transform 1 0 49036 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_529
timestamp 1666464484
transform 1 0 49772 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_537
timestamp 1666464484
transform 1 0 50508 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_545
timestamp 1666464484
transform 1 0 51244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_553
timestamp 1666464484
transform 1 0 51980 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_557
timestamp 1666464484
transform 1 0 52348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1666464484
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_561
timestamp 1666464484
transform 1 0 52716 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_569
timestamp 1666464484
transform 1 0 53452 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_577
timestamp 1666464484
transform 1 0 54188 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_585
timestamp 1666464484
transform 1 0 54924 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_593
timestamp 1666464484
transform 1 0 55660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_53_601
timestamp 1666464484
transform 1 0 56396 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_609
timestamp 1666464484
transform 1 0 57132 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_613
timestamp 1666464484
transform 1 0 57500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1666464484
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_617
timestamp 1666464484
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_3
timestamp 1666464484
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_11
timestamp 1666464484
transform 1 0 2116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_19
timestamp 1666464484
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1666464484
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_29
timestamp 1666464484
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_37
timestamp 1666464484
transform 1 0 4508 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_45
timestamp 1666464484
transform 1 0 5244 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_53
timestamp 1666464484
transform 1 0 5980 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_61
timestamp 1666464484
transform 1 0 6716 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_69
timestamp 1666464484
transform 1 0 7452 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_77
timestamp 1666464484
transform 1 0 8188 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_81
timestamp 1666464484
transform 1 0 8556 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1666464484
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_85
timestamp 1666464484
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_93
timestamp 1666464484
transform 1 0 9660 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_101
timestamp 1666464484
transform 1 0 10396 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_109
timestamp 1666464484
transform 1 0 11132 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_117
timestamp 1666464484
transform 1 0 11868 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_125
timestamp 1666464484
transform 1 0 12604 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_133
timestamp 1666464484
transform 1 0 13340 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_137
timestamp 1666464484
transform 1 0 13708 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1666464484
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_141
timestamp 1666464484
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_149
timestamp 1666464484
transform 1 0 14812 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_157
timestamp 1666464484
transform 1 0 15548 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_165
timestamp 1666464484
transform 1 0 16284 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_173
timestamp 1666464484
transform 1 0 17020 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_181
timestamp 1666464484
transform 1 0 17756 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_189
timestamp 1666464484
transform 1 0 18492 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_193
timestamp 1666464484
transform 1 0 18860 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1666464484
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_197
timestamp 1666464484
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_205
timestamp 1666464484
transform 1 0 19964 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_213
timestamp 1666464484
transform 1 0 20700 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_221
timestamp 1666464484
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_229
timestamp 1666464484
transform 1 0 22172 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_237
timestamp 1666464484
transform 1 0 22908 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_245
timestamp 1666464484
transform 1 0 23644 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_249
timestamp 1666464484
transform 1 0 24012 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1666464484
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_253
timestamp 1666464484
transform 1 0 24380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_261
timestamp 1666464484
transform 1 0 25116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_269
timestamp 1666464484
transform 1 0 25852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_277
timestamp 1666464484
transform 1 0 26588 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_285
timestamp 1666464484
transform 1 0 27324 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_293
timestamp 1666464484
transform 1 0 28060 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_301
timestamp 1666464484
transform 1 0 28796 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_305
timestamp 1666464484
transform 1 0 29164 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1666464484
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_309
timestamp 1666464484
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_317
timestamp 1666464484
transform 1 0 30268 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_325
timestamp 1666464484
transform 1 0 31004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_333
timestamp 1666464484
transform 1 0 31740 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_341
timestamp 1666464484
transform 1 0 32476 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_349
timestamp 1666464484
transform 1 0 33212 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_357
timestamp 1666464484
transform 1 0 33948 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_361
timestamp 1666464484
transform 1 0 34316 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1666464484
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_365
timestamp 1666464484
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_373
timestamp 1666464484
transform 1 0 35420 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_381
timestamp 1666464484
transform 1 0 36156 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_389
timestamp 1666464484
transform 1 0 36892 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_397
timestamp 1666464484
transform 1 0 37628 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_405
timestamp 1666464484
transform 1 0 38364 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_413
timestamp 1666464484
transform 1 0 39100 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_417
timestamp 1666464484
transform 1 0 39468 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1666464484
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_421
timestamp 1666464484
transform 1 0 39836 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_429
timestamp 1666464484
transform 1 0 40572 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_437
timestamp 1666464484
transform 1 0 41308 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_445
timestamp 1666464484
transform 1 0 42044 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_453
timestamp 1666464484
transform 1 0 42780 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_461
timestamp 1666464484
transform 1 0 43516 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_469
timestamp 1666464484
transform 1 0 44252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_473
timestamp 1666464484
transform 1 0 44620 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1666464484
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_477
timestamp 1666464484
transform 1 0 44988 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_485
timestamp 1666464484
transform 1 0 45724 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_493
timestamp 1666464484
transform 1 0 46460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_501
timestamp 1666464484
transform 1 0 47196 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_509
timestamp 1666464484
transform 1 0 47932 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_517
timestamp 1666464484
transform 1 0 48668 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_525
timestamp 1666464484
transform 1 0 49404 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_529
timestamp 1666464484
transform 1 0 49772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1666464484
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_533
timestamp 1666464484
transform 1 0 50140 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_541
timestamp 1666464484
transform 1 0 50876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_549
timestamp 1666464484
transform 1 0 51612 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_557
timestamp 1666464484
transform 1 0 52348 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_565
timestamp 1666464484
transform 1 0 53084 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_573
timestamp 1666464484
transform 1 0 53820 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_581
timestamp 1666464484
transform 1 0 54556 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_585
timestamp 1666464484
transform 1 0 54924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1666464484
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_589
timestamp 1666464484
transform 1 0 55292 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_597
timestamp 1666464484
transform 1 0 56028 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_605
timestamp 1666464484
transform 1 0 56764 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_54_613
timestamp 1666464484
transform 1 0 57500 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_621
timestamp 1666464484
transform 1 0 58236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_55_3
timestamp 1666464484
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_11
timestamp 1666464484
transform 1 0 2116 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_19
timestamp 1666464484
transform 1 0 2852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_27
timestamp 1666464484
transform 1 0 3588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_35
timestamp 1666464484
transform 1 0 4324 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_43
timestamp 1666464484
transform 1 0 5060 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_51
timestamp 1666464484
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1666464484
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_57
timestamp 1666464484
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_65
timestamp 1666464484
transform 1 0 7084 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_73
timestamp 1666464484
transform 1 0 7820 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_81
timestamp 1666464484
transform 1 0 8556 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_89
timestamp 1666464484
transform 1 0 9292 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_97
timestamp 1666464484
transform 1 0 10028 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_105
timestamp 1666464484
transform 1 0 10764 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_109
timestamp 1666464484
transform 1 0 11132 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1666464484
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_113
timestamp 1666464484
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_121
timestamp 1666464484
transform 1 0 12236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_129
timestamp 1666464484
transform 1 0 12972 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_137
timestamp 1666464484
transform 1 0 13708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_145
timestamp 1666464484
transform 1 0 14444 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_153
timestamp 1666464484
transform 1 0 15180 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_161
timestamp 1666464484
transform 1 0 15916 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_165
timestamp 1666464484
transform 1 0 16284 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1666464484
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_169
timestamp 1666464484
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_177
timestamp 1666464484
transform 1 0 17388 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_185
timestamp 1666464484
transform 1 0 18124 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_193
timestamp 1666464484
transform 1 0 18860 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_201
timestamp 1666464484
transform 1 0 19596 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_209
timestamp 1666464484
transform 1 0 20332 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_217
timestamp 1666464484
transform 1 0 21068 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_221
timestamp 1666464484
transform 1 0 21436 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1666464484
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_225
timestamp 1666464484
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_233
timestamp 1666464484
transform 1 0 22540 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_241
timestamp 1666464484
transform 1 0 23276 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_249
timestamp 1666464484
transform 1 0 24012 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_257
timestamp 1666464484
transform 1 0 24748 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_265
timestamp 1666464484
transform 1 0 25484 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_273
timestamp 1666464484
transform 1 0 26220 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_277
timestamp 1666464484
transform 1 0 26588 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1666464484
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_281
timestamp 1666464484
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_289
timestamp 1666464484
transform 1 0 27692 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_297
timestamp 1666464484
transform 1 0 28428 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_305
timestamp 1666464484
transform 1 0 29164 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_313
timestamp 1666464484
transform 1 0 29900 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_321
timestamp 1666464484
transform 1 0 30636 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_329
timestamp 1666464484
transform 1 0 31372 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_333
timestamp 1666464484
transform 1 0 31740 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1666464484
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_337
timestamp 1666464484
transform 1 0 32108 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_345
timestamp 1666464484
transform 1 0 32844 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_353
timestamp 1666464484
transform 1 0 33580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_361
timestamp 1666464484
transform 1 0 34316 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_369
timestamp 1666464484
transform 1 0 35052 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_377
timestamp 1666464484
transform 1 0 35788 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_385
timestamp 1666464484
transform 1 0 36524 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_389
timestamp 1666464484
transform 1 0 36892 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1666464484
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_393
timestamp 1666464484
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_401
timestamp 1666464484
transform 1 0 37996 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_409
timestamp 1666464484
transform 1 0 38732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_417
timestamp 1666464484
transform 1 0 39468 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_425
timestamp 1666464484
transform 1 0 40204 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_433
timestamp 1666464484
transform 1 0 40940 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_441
timestamp 1666464484
transform 1 0 41676 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_445
timestamp 1666464484
transform 1 0 42044 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1666464484
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_449
timestamp 1666464484
transform 1 0 42412 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_457
timestamp 1666464484
transform 1 0 43148 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_465
timestamp 1666464484
transform 1 0 43884 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_473
timestamp 1666464484
transform 1 0 44620 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_481
timestamp 1666464484
transform 1 0 45356 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_489
timestamp 1666464484
transform 1 0 46092 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_497
timestamp 1666464484
transform 1 0 46828 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_501
timestamp 1666464484
transform 1 0 47196 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1666464484
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_505
timestamp 1666464484
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_513
timestamp 1666464484
transform 1 0 48300 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_521
timestamp 1666464484
transform 1 0 49036 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_529
timestamp 1666464484
transform 1 0 49772 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_537
timestamp 1666464484
transform 1 0 50508 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_545
timestamp 1666464484
transform 1 0 51244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_553
timestamp 1666464484
transform 1 0 51980 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_557
timestamp 1666464484
transform 1 0 52348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1666464484
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_561
timestamp 1666464484
transform 1 0 52716 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_569
timestamp 1666464484
transform 1 0 53452 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_577
timestamp 1666464484
transform 1 0 54188 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_585
timestamp 1666464484
transform 1 0 54924 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_593
timestamp 1666464484
transform 1 0 55660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_601
timestamp 1666464484
transform 1 0 56396 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_609
timestamp 1666464484
transform 1 0 57132 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_613
timestamp 1666464484
transform 1 0 57500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1666464484
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_617
timestamp 1666464484
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_3
timestamp 1666464484
transform 1 0 1380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_11
timestamp 1666464484
transform 1 0 2116 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_19
timestamp 1666464484
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1666464484
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_29
timestamp 1666464484
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_37
timestamp 1666464484
transform 1 0 4508 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_45
timestamp 1666464484
transform 1 0 5244 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_53
timestamp 1666464484
transform 1 0 5980 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_61
timestamp 1666464484
transform 1 0 6716 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_69
timestamp 1666464484
transform 1 0 7452 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_77
timestamp 1666464484
transform 1 0 8188 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_81
timestamp 1666464484
transform 1 0 8556 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1666464484
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_85
timestamp 1666464484
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_93
timestamp 1666464484
transform 1 0 9660 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_101
timestamp 1666464484
transform 1 0 10396 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_109
timestamp 1666464484
transform 1 0 11132 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_117
timestamp 1666464484
transform 1 0 11868 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_125
timestamp 1666464484
transform 1 0 12604 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_133
timestamp 1666464484
transform 1 0 13340 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_137
timestamp 1666464484
transform 1 0 13708 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1666464484
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_141
timestamp 1666464484
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_149
timestamp 1666464484
transform 1 0 14812 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_157
timestamp 1666464484
transform 1 0 15548 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_165
timestamp 1666464484
transform 1 0 16284 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_173
timestamp 1666464484
transform 1 0 17020 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_181
timestamp 1666464484
transform 1 0 17756 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_189
timestamp 1666464484
transform 1 0 18492 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_193
timestamp 1666464484
transform 1 0 18860 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1666464484
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_197
timestamp 1666464484
transform 1 0 19228 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_205
timestamp 1666464484
transform 1 0 19964 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_213
timestamp 1666464484
transform 1 0 20700 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_221
timestamp 1666464484
transform 1 0 21436 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_229
timestamp 1666464484
transform 1 0 22172 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_237
timestamp 1666464484
transform 1 0 22908 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_245
timestamp 1666464484
transform 1 0 23644 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_249
timestamp 1666464484
transform 1 0 24012 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1666464484
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_253
timestamp 1666464484
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_261
timestamp 1666464484
transform 1 0 25116 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_269
timestamp 1666464484
transform 1 0 25852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_277
timestamp 1666464484
transform 1 0 26588 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_285
timestamp 1666464484
transform 1 0 27324 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_293
timestamp 1666464484
transform 1 0 28060 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_301
timestamp 1666464484
transform 1 0 28796 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_305
timestamp 1666464484
transform 1 0 29164 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1666464484
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_309
timestamp 1666464484
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_317
timestamp 1666464484
transform 1 0 30268 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_325
timestamp 1666464484
transform 1 0 31004 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_333
timestamp 1666464484
transform 1 0 31740 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_341
timestamp 1666464484
transform 1 0 32476 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_349
timestamp 1666464484
transform 1 0 33212 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_357
timestamp 1666464484
transform 1 0 33948 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_361
timestamp 1666464484
transform 1 0 34316 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1666464484
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_365
timestamp 1666464484
transform 1 0 34684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_373
timestamp 1666464484
transform 1 0 35420 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_381
timestamp 1666464484
transform 1 0 36156 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_389
timestamp 1666464484
transform 1 0 36892 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_397
timestamp 1666464484
transform 1 0 37628 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_405
timestamp 1666464484
transform 1 0 38364 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_413
timestamp 1666464484
transform 1 0 39100 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_417
timestamp 1666464484
transform 1 0 39468 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1666464484
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_421
timestamp 1666464484
transform 1 0 39836 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_429
timestamp 1666464484
transform 1 0 40572 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_437
timestamp 1666464484
transform 1 0 41308 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_445
timestamp 1666464484
transform 1 0 42044 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_453
timestamp 1666464484
transform 1 0 42780 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_461
timestamp 1666464484
transform 1 0 43516 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_469
timestamp 1666464484
transform 1 0 44252 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_473
timestamp 1666464484
transform 1 0 44620 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1666464484
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_477
timestamp 1666464484
transform 1 0 44988 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_485
timestamp 1666464484
transform 1 0 45724 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_493
timestamp 1666464484
transform 1 0 46460 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_501
timestamp 1666464484
transform 1 0 47196 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_509
timestamp 1666464484
transform 1 0 47932 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_517
timestamp 1666464484
transform 1 0 48668 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_525
timestamp 1666464484
transform 1 0 49404 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_529
timestamp 1666464484
transform 1 0 49772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1666464484
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_533
timestamp 1666464484
transform 1 0 50140 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_541
timestamp 1666464484
transform 1 0 50876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_549
timestamp 1666464484
transform 1 0 51612 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_557
timestamp 1666464484
transform 1 0 52348 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_565
timestamp 1666464484
transform 1 0 53084 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_573
timestamp 1666464484
transform 1 0 53820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_581
timestamp 1666464484
transform 1 0 54556 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_585
timestamp 1666464484
transform 1 0 54924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1666464484
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_56_589
timestamp 1666464484
transform 1 0 55292 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_597
timestamp 1666464484
transform 1 0 56028 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_605
timestamp 1666464484
transform 1 0 56764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_56_613
timestamp 1666464484
transform 1 0 57500 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_621
timestamp 1666464484
transform 1 0 58236 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_57_3
timestamp 1666464484
transform 1 0 1380 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_11
timestamp 1666464484
transform 1 0 2116 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_19
timestamp 1666464484
transform 1 0 2852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_27
timestamp 1666464484
transform 1 0 3588 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_35
timestamp 1666464484
transform 1 0 4324 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_43
timestamp 1666464484
transform 1 0 5060 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_51
timestamp 1666464484
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1666464484
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_57
timestamp 1666464484
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_65
timestamp 1666464484
transform 1 0 7084 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_73
timestamp 1666464484
transform 1 0 7820 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_81
timestamp 1666464484
transform 1 0 8556 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_89
timestamp 1666464484
transform 1 0 9292 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_97
timestamp 1666464484
transform 1 0 10028 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_105
timestamp 1666464484
transform 1 0 10764 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_109
timestamp 1666464484
transform 1 0 11132 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1666464484
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_113
timestamp 1666464484
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_121
timestamp 1666464484
transform 1 0 12236 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_129
timestamp 1666464484
transform 1 0 12972 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_137
timestamp 1666464484
transform 1 0 13708 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_145
timestamp 1666464484
transform 1 0 14444 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_153
timestamp 1666464484
transform 1 0 15180 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_161
timestamp 1666464484
transform 1 0 15916 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_165
timestamp 1666464484
transform 1 0 16284 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1666464484
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_169
timestamp 1666464484
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_177
timestamp 1666464484
transform 1 0 17388 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_185
timestamp 1666464484
transform 1 0 18124 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_193
timestamp 1666464484
transform 1 0 18860 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_201
timestamp 1666464484
transform 1 0 19596 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_209
timestamp 1666464484
transform 1 0 20332 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_217
timestamp 1666464484
transform 1 0 21068 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_221
timestamp 1666464484
transform 1 0 21436 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1666464484
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_225
timestamp 1666464484
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_233
timestamp 1666464484
transform 1 0 22540 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_241
timestamp 1666464484
transform 1 0 23276 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_249
timestamp 1666464484
transform 1 0 24012 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_257
timestamp 1666464484
transform 1 0 24748 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_265
timestamp 1666464484
transform 1 0 25484 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_273
timestamp 1666464484
transform 1 0 26220 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_277
timestamp 1666464484
transform 1 0 26588 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1666464484
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_281
timestamp 1666464484
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_289
timestamp 1666464484
transform 1 0 27692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_297
timestamp 1666464484
transform 1 0 28428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_305
timestamp 1666464484
transform 1 0 29164 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_313
timestamp 1666464484
transform 1 0 29900 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_321
timestamp 1666464484
transform 1 0 30636 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_329
timestamp 1666464484
transform 1 0 31372 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_333
timestamp 1666464484
transform 1 0 31740 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1666464484
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_337
timestamp 1666464484
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_345
timestamp 1666464484
transform 1 0 32844 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_353
timestamp 1666464484
transform 1 0 33580 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_361
timestamp 1666464484
transform 1 0 34316 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_369
timestamp 1666464484
transform 1 0 35052 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_377
timestamp 1666464484
transform 1 0 35788 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_385
timestamp 1666464484
transform 1 0 36524 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_389
timestamp 1666464484
transform 1 0 36892 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1666464484
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_393
timestamp 1666464484
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_401
timestamp 1666464484
transform 1 0 37996 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_409
timestamp 1666464484
transform 1 0 38732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_417
timestamp 1666464484
transform 1 0 39468 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_425
timestamp 1666464484
transform 1 0 40204 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_433
timestamp 1666464484
transform 1 0 40940 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_441
timestamp 1666464484
transform 1 0 41676 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_445
timestamp 1666464484
transform 1 0 42044 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1666464484
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_449
timestamp 1666464484
transform 1 0 42412 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_457
timestamp 1666464484
transform 1 0 43148 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_465
timestamp 1666464484
transform 1 0 43884 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_473
timestamp 1666464484
transform 1 0 44620 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_481
timestamp 1666464484
transform 1 0 45356 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_489
timestamp 1666464484
transform 1 0 46092 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_497
timestamp 1666464484
transform 1 0 46828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_501
timestamp 1666464484
transform 1 0 47196 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1666464484
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_505
timestamp 1666464484
transform 1 0 47564 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_513
timestamp 1666464484
transform 1 0 48300 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_521
timestamp 1666464484
transform 1 0 49036 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_529
timestamp 1666464484
transform 1 0 49772 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_537
timestamp 1666464484
transform 1 0 50508 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_545
timestamp 1666464484
transform 1 0 51244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_553
timestamp 1666464484
transform 1 0 51980 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_557
timestamp 1666464484
transform 1 0 52348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1666464484
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_561
timestamp 1666464484
transform 1 0 52716 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_569
timestamp 1666464484
transform 1 0 53452 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_577
timestamp 1666464484
transform 1 0 54188 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_585
timestamp 1666464484
transform 1 0 54924 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_593
timestamp 1666464484
transform 1 0 55660 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_57_601
timestamp 1666464484
transform 1 0 56396 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_609
timestamp 1666464484
transform 1 0 57132 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_613
timestamp 1666464484
transform 1 0 57500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1666464484
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_57_617
timestamp 1666464484
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_3
timestamp 1666464484
transform 1 0 1380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_11
timestamp 1666464484
transform 1 0 2116 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_19
timestamp 1666464484
transform 1 0 2852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1666464484
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_29
timestamp 1666464484
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_37
timestamp 1666464484
transform 1 0 4508 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_45
timestamp 1666464484
transform 1 0 5244 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_53
timestamp 1666464484
transform 1 0 5980 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_61
timestamp 1666464484
transform 1 0 6716 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_69
timestamp 1666464484
transform 1 0 7452 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_77
timestamp 1666464484
transform 1 0 8188 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_81
timestamp 1666464484
transform 1 0 8556 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1666464484
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_85
timestamp 1666464484
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_93
timestamp 1666464484
transform 1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_101
timestamp 1666464484
transform 1 0 10396 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_109
timestamp 1666464484
transform 1 0 11132 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_117
timestamp 1666464484
transform 1 0 11868 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_125
timestamp 1666464484
transform 1 0 12604 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_133
timestamp 1666464484
transform 1 0 13340 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_137
timestamp 1666464484
transform 1 0 13708 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1666464484
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_141
timestamp 1666464484
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_149
timestamp 1666464484
transform 1 0 14812 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_157
timestamp 1666464484
transform 1 0 15548 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_165
timestamp 1666464484
transform 1 0 16284 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_173
timestamp 1666464484
transform 1 0 17020 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_181
timestamp 1666464484
transform 1 0 17756 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_189
timestamp 1666464484
transform 1 0 18492 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_193
timestamp 1666464484
transform 1 0 18860 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1666464484
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_197
timestamp 1666464484
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_205
timestamp 1666464484
transform 1 0 19964 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_213
timestamp 1666464484
transform 1 0 20700 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_221
timestamp 1666464484
transform 1 0 21436 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_229
timestamp 1666464484
transform 1 0 22172 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_237
timestamp 1666464484
transform 1 0 22908 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_245
timestamp 1666464484
transform 1 0 23644 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_249
timestamp 1666464484
transform 1 0 24012 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1666464484
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_253
timestamp 1666464484
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_261
timestamp 1666464484
transform 1 0 25116 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_269
timestamp 1666464484
transform 1 0 25852 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_277
timestamp 1666464484
transform 1 0 26588 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_285
timestamp 1666464484
transform 1 0 27324 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_293
timestamp 1666464484
transform 1 0 28060 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_301
timestamp 1666464484
transform 1 0 28796 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_305
timestamp 1666464484
transform 1 0 29164 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1666464484
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_309
timestamp 1666464484
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_317
timestamp 1666464484
transform 1 0 30268 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_325
timestamp 1666464484
transform 1 0 31004 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_333
timestamp 1666464484
transform 1 0 31740 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_341
timestamp 1666464484
transform 1 0 32476 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_349
timestamp 1666464484
transform 1 0 33212 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_357
timestamp 1666464484
transform 1 0 33948 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_361
timestamp 1666464484
transform 1 0 34316 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1666464484
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_365
timestamp 1666464484
transform 1 0 34684 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_373
timestamp 1666464484
transform 1 0 35420 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_381
timestamp 1666464484
transform 1 0 36156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_389
timestamp 1666464484
transform 1 0 36892 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_397
timestamp 1666464484
transform 1 0 37628 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_405
timestamp 1666464484
transform 1 0 38364 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_413
timestamp 1666464484
transform 1 0 39100 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_417
timestamp 1666464484
transform 1 0 39468 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1666464484
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_421
timestamp 1666464484
transform 1 0 39836 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_429
timestamp 1666464484
transform 1 0 40572 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_437
timestamp 1666464484
transform 1 0 41308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_445
timestamp 1666464484
transform 1 0 42044 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_453
timestamp 1666464484
transform 1 0 42780 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_461
timestamp 1666464484
transform 1 0 43516 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_469
timestamp 1666464484
transform 1 0 44252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_473
timestamp 1666464484
transform 1 0 44620 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1666464484
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_477
timestamp 1666464484
transform 1 0 44988 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_485
timestamp 1666464484
transform 1 0 45724 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_493
timestamp 1666464484
transform 1 0 46460 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_501
timestamp 1666464484
transform 1 0 47196 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_509
timestamp 1666464484
transform 1 0 47932 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_517
timestamp 1666464484
transform 1 0 48668 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_525
timestamp 1666464484
transform 1 0 49404 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_529
timestamp 1666464484
transform 1 0 49772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1666464484
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_533
timestamp 1666464484
transform 1 0 50140 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_541
timestamp 1666464484
transform 1 0 50876 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_549
timestamp 1666464484
transform 1 0 51612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_557
timestamp 1666464484
transform 1 0 52348 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_565
timestamp 1666464484
transform 1 0 53084 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_573
timestamp 1666464484
transform 1 0 53820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_581
timestamp 1666464484
transform 1 0 54556 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_585
timestamp 1666464484
transform 1 0 54924 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1666464484
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_589
timestamp 1666464484
transform 1 0 55292 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_597
timestamp 1666464484
transform 1 0 56028 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_605
timestamp 1666464484
transform 1 0 56764 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_58_613
timestamp 1666464484
transform 1 0 57500 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_621
timestamp 1666464484
transform 1 0 58236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_59_3
timestamp 1666464484
transform 1 0 1380 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_11
timestamp 1666464484
transform 1 0 2116 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_19
timestamp 1666464484
transform 1 0 2852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_27
timestamp 1666464484
transform 1 0 3588 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_35
timestamp 1666464484
transform 1 0 4324 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_43
timestamp 1666464484
transform 1 0 5060 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_51
timestamp 1666464484
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1666464484
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_57
timestamp 1666464484
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_65
timestamp 1666464484
transform 1 0 7084 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_73
timestamp 1666464484
transform 1 0 7820 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_81
timestamp 1666464484
transform 1 0 8556 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_89
timestamp 1666464484
transform 1 0 9292 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_97
timestamp 1666464484
transform 1 0 10028 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_105
timestamp 1666464484
transform 1 0 10764 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_109
timestamp 1666464484
transform 1 0 11132 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1666464484
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_113
timestamp 1666464484
transform 1 0 11500 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_121
timestamp 1666464484
transform 1 0 12236 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_129
timestamp 1666464484
transform 1 0 12972 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_137
timestamp 1666464484
transform 1 0 13708 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_145
timestamp 1666464484
transform 1 0 14444 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_153
timestamp 1666464484
transform 1 0 15180 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_161
timestamp 1666464484
transform 1 0 15916 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_165
timestamp 1666464484
transform 1 0 16284 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1666464484
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_169
timestamp 1666464484
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_177
timestamp 1666464484
transform 1 0 17388 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_185
timestamp 1666464484
transform 1 0 18124 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_193
timestamp 1666464484
transform 1 0 18860 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_201
timestamp 1666464484
transform 1 0 19596 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_209
timestamp 1666464484
transform 1 0 20332 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_217
timestamp 1666464484
transform 1 0 21068 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_221
timestamp 1666464484
transform 1 0 21436 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1666464484
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_225
timestamp 1666464484
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_233
timestamp 1666464484
transform 1 0 22540 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_241
timestamp 1666464484
transform 1 0 23276 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_249
timestamp 1666464484
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_257
timestamp 1666464484
transform 1 0 24748 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_265
timestamp 1666464484
transform 1 0 25484 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_273
timestamp 1666464484
transform 1 0 26220 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_277
timestamp 1666464484
transform 1 0 26588 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1666464484
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_281
timestamp 1666464484
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_289
timestamp 1666464484
transform 1 0 27692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_297
timestamp 1666464484
transform 1 0 28428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_305
timestamp 1666464484
transform 1 0 29164 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_313
timestamp 1666464484
transform 1 0 29900 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_321
timestamp 1666464484
transform 1 0 30636 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_329
timestamp 1666464484
transform 1 0 31372 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_333
timestamp 1666464484
transform 1 0 31740 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1666464484
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_337
timestamp 1666464484
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_345
timestamp 1666464484
transform 1 0 32844 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_353
timestamp 1666464484
transform 1 0 33580 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_361
timestamp 1666464484
transform 1 0 34316 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_369
timestamp 1666464484
transform 1 0 35052 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_377
timestamp 1666464484
transform 1 0 35788 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_385
timestamp 1666464484
transform 1 0 36524 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_389
timestamp 1666464484
transform 1 0 36892 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1666464484
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_393
timestamp 1666464484
transform 1 0 37260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_401
timestamp 1666464484
transform 1 0 37996 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_409
timestamp 1666464484
transform 1 0 38732 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_417
timestamp 1666464484
transform 1 0 39468 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_425
timestamp 1666464484
transform 1 0 40204 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_433
timestamp 1666464484
transform 1 0 40940 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_441
timestamp 1666464484
transform 1 0 41676 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_445
timestamp 1666464484
transform 1 0 42044 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1666464484
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_449
timestamp 1666464484
transform 1 0 42412 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_457
timestamp 1666464484
transform 1 0 43148 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_465
timestamp 1666464484
transform 1 0 43884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_473
timestamp 1666464484
transform 1 0 44620 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_481
timestamp 1666464484
transform 1 0 45356 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_489
timestamp 1666464484
transform 1 0 46092 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_497
timestamp 1666464484
transform 1 0 46828 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_501
timestamp 1666464484
transform 1 0 47196 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1666464484
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_505
timestamp 1666464484
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_513
timestamp 1666464484
transform 1 0 48300 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_521
timestamp 1666464484
transform 1 0 49036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_529
timestamp 1666464484
transform 1 0 49772 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_537
timestamp 1666464484
transform 1 0 50508 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_545
timestamp 1666464484
transform 1 0 51244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_553
timestamp 1666464484
transform 1 0 51980 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_557
timestamp 1666464484
transform 1 0 52348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1666464484
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_561
timestamp 1666464484
transform 1 0 52716 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_569
timestamp 1666464484
transform 1 0 53452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_577
timestamp 1666464484
transform 1 0 54188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_585
timestamp 1666464484
transform 1 0 54924 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_593
timestamp 1666464484
transform 1 0 55660 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_59_601
timestamp 1666464484
transform 1 0 56396 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_609
timestamp 1666464484
transform 1 0 57132 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_613
timestamp 1666464484
transform 1 0 57500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1666464484
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_59_617
timestamp 1666464484
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_3
timestamp 1666464484
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_11
timestamp 1666464484
transform 1 0 2116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_19
timestamp 1666464484
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1666464484
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_29
timestamp 1666464484
transform 1 0 3772 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_37
timestamp 1666464484
transform 1 0 4508 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_45
timestamp 1666464484
transform 1 0 5244 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_53
timestamp 1666464484
transform 1 0 5980 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_61
timestamp 1666464484
transform 1 0 6716 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_69
timestamp 1666464484
transform 1 0 7452 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_77
timestamp 1666464484
transform 1 0 8188 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_81
timestamp 1666464484
transform 1 0 8556 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1666464484
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_85
timestamp 1666464484
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_93
timestamp 1666464484
transform 1 0 9660 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_101
timestamp 1666464484
transform 1 0 10396 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_109
timestamp 1666464484
transform 1 0 11132 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_117
timestamp 1666464484
transform 1 0 11868 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_125
timestamp 1666464484
transform 1 0 12604 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_133
timestamp 1666464484
transform 1 0 13340 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_137
timestamp 1666464484
transform 1 0 13708 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1666464484
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_141
timestamp 1666464484
transform 1 0 14076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_149
timestamp 1666464484
transform 1 0 14812 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_157
timestamp 1666464484
transform 1 0 15548 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_165
timestamp 1666464484
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_173
timestamp 1666464484
transform 1 0 17020 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_181
timestamp 1666464484
transform 1 0 17756 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_189
timestamp 1666464484
transform 1 0 18492 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_193
timestamp 1666464484
transform 1 0 18860 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1666464484
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_197
timestamp 1666464484
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_205
timestamp 1666464484
transform 1 0 19964 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_213
timestamp 1666464484
transform 1 0 20700 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_221
timestamp 1666464484
transform 1 0 21436 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_229
timestamp 1666464484
transform 1 0 22172 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_237
timestamp 1666464484
transform 1 0 22908 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_245
timestamp 1666464484
transform 1 0 23644 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_249
timestamp 1666464484
transform 1 0 24012 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1666464484
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_253
timestamp 1666464484
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_261
timestamp 1666464484
transform 1 0 25116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_269
timestamp 1666464484
transform 1 0 25852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_277
timestamp 1666464484
transform 1 0 26588 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_285
timestamp 1666464484
transform 1 0 27324 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_293
timestamp 1666464484
transform 1 0 28060 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_301
timestamp 1666464484
transform 1 0 28796 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_305
timestamp 1666464484
transform 1 0 29164 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1666464484
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_309
timestamp 1666464484
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_317
timestamp 1666464484
transform 1 0 30268 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_325
timestamp 1666464484
transform 1 0 31004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_333
timestamp 1666464484
transform 1 0 31740 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_341
timestamp 1666464484
transform 1 0 32476 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_349
timestamp 1666464484
transform 1 0 33212 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_357
timestamp 1666464484
transform 1 0 33948 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_361
timestamp 1666464484
transform 1 0 34316 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1666464484
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_365
timestamp 1666464484
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_373
timestamp 1666464484
transform 1 0 35420 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_381
timestamp 1666464484
transform 1 0 36156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_389
timestamp 1666464484
transform 1 0 36892 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_397
timestamp 1666464484
transform 1 0 37628 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_405
timestamp 1666464484
transform 1 0 38364 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_413
timestamp 1666464484
transform 1 0 39100 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_417
timestamp 1666464484
transform 1 0 39468 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1666464484
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_421
timestamp 1666464484
transform 1 0 39836 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_429
timestamp 1666464484
transform 1 0 40572 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_437
timestamp 1666464484
transform 1 0 41308 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_445
timestamp 1666464484
transform 1 0 42044 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_453
timestamp 1666464484
transform 1 0 42780 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_461
timestamp 1666464484
transform 1 0 43516 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_469
timestamp 1666464484
transform 1 0 44252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_473
timestamp 1666464484
transform 1 0 44620 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1666464484
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_477
timestamp 1666464484
transform 1 0 44988 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_485
timestamp 1666464484
transform 1 0 45724 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_493
timestamp 1666464484
transform 1 0 46460 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_501
timestamp 1666464484
transform 1 0 47196 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_509
timestamp 1666464484
transform 1 0 47932 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_517
timestamp 1666464484
transform 1 0 48668 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_525
timestamp 1666464484
transform 1 0 49404 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_529
timestamp 1666464484
transform 1 0 49772 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1666464484
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_533
timestamp 1666464484
transform 1 0 50140 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_541
timestamp 1666464484
transform 1 0 50876 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_549
timestamp 1666464484
transform 1 0 51612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_557
timestamp 1666464484
transform 1 0 52348 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_565
timestamp 1666464484
transform 1 0 53084 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_573
timestamp 1666464484
transform 1 0 53820 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_581
timestamp 1666464484
transform 1 0 54556 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_585
timestamp 1666464484
transform 1 0 54924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1666464484
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_589
timestamp 1666464484
transform 1 0 55292 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_597
timestamp 1666464484
transform 1 0 56028 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_605
timestamp 1666464484
transform 1 0 56764 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_613
timestamp 1666464484
transform 1 0 57500 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_621
timestamp 1666464484
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_61_3
timestamp 1666464484
transform 1 0 1380 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_11
timestamp 1666464484
transform 1 0 2116 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_19
timestamp 1666464484
transform 1 0 2852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_27
timestamp 1666464484
transform 1 0 3588 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_35
timestamp 1666464484
transform 1 0 4324 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_43
timestamp 1666464484
transform 1 0 5060 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_51
timestamp 1666464484
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1666464484
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_57
timestamp 1666464484
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_65
timestamp 1666464484
transform 1 0 7084 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_73
timestamp 1666464484
transform 1 0 7820 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_81
timestamp 1666464484
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_89
timestamp 1666464484
transform 1 0 9292 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_97
timestamp 1666464484
transform 1 0 10028 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_105
timestamp 1666464484
transform 1 0 10764 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_109
timestamp 1666464484
transform 1 0 11132 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1666464484
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_113
timestamp 1666464484
transform 1 0 11500 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_121
timestamp 1666464484
transform 1 0 12236 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_129
timestamp 1666464484
transform 1 0 12972 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_137
timestamp 1666464484
transform 1 0 13708 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_145
timestamp 1666464484
transform 1 0 14444 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_153
timestamp 1666464484
transform 1 0 15180 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_161
timestamp 1666464484
transform 1 0 15916 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_165
timestamp 1666464484
transform 1 0 16284 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1666464484
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_169
timestamp 1666464484
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_177
timestamp 1666464484
transform 1 0 17388 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_185
timestamp 1666464484
transform 1 0 18124 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_193
timestamp 1666464484
transform 1 0 18860 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_201
timestamp 1666464484
transform 1 0 19596 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_209
timestamp 1666464484
transform 1 0 20332 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_217
timestamp 1666464484
transform 1 0 21068 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_221
timestamp 1666464484
transform 1 0 21436 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1666464484
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_225
timestamp 1666464484
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_233
timestamp 1666464484
transform 1 0 22540 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_241
timestamp 1666464484
transform 1 0 23276 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_249
timestamp 1666464484
transform 1 0 24012 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_257
timestamp 1666464484
transform 1 0 24748 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_265
timestamp 1666464484
transform 1 0 25484 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_273
timestamp 1666464484
transform 1 0 26220 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_277
timestamp 1666464484
transform 1 0 26588 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1666464484
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_281
timestamp 1666464484
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_289
timestamp 1666464484
transform 1 0 27692 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_297
timestamp 1666464484
transform 1 0 28428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_305
timestamp 1666464484
transform 1 0 29164 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_313
timestamp 1666464484
transform 1 0 29900 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_321
timestamp 1666464484
transform 1 0 30636 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_329
timestamp 1666464484
transform 1 0 31372 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_333
timestamp 1666464484
transform 1 0 31740 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1666464484
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_337
timestamp 1666464484
transform 1 0 32108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_345
timestamp 1666464484
transform 1 0 32844 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_353
timestamp 1666464484
transform 1 0 33580 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_361
timestamp 1666464484
transform 1 0 34316 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_369
timestamp 1666464484
transform 1 0 35052 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_377
timestamp 1666464484
transform 1 0 35788 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_385
timestamp 1666464484
transform 1 0 36524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_389
timestamp 1666464484
transform 1 0 36892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1666464484
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_393
timestamp 1666464484
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_401
timestamp 1666464484
transform 1 0 37996 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_409
timestamp 1666464484
transform 1 0 38732 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_417
timestamp 1666464484
transform 1 0 39468 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_425
timestamp 1666464484
transform 1 0 40204 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_433
timestamp 1666464484
transform 1 0 40940 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_441
timestamp 1666464484
transform 1 0 41676 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_445
timestamp 1666464484
transform 1 0 42044 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1666464484
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_449
timestamp 1666464484
transform 1 0 42412 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_457
timestamp 1666464484
transform 1 0 43148 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_465
timestamp 1666464484
transform 1 0 43884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_473
timestamp 1666464484
transform 1 0 44620 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_481
timestamp 1666464484
transform 1 0 45356 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_489
timestamp 1666464484
transform 1 0 46092 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_497
timestamp 1666464484
transform 1 0 46828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_501
timestamp 1666464484
transform 1 0 47196 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1666464484
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_505
timestamp 1666464484
transform 1 0 47564 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_513
timestamp 1666464484
transform 1 0 48300 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_521
timestamp 1666464484
transform 1 0 49036 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_529
timestamp 1666464484
transform 1 0 49772 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_537
timestamp 1666464484
transform 1 0 50508 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_545
timestamp 1666464484
transform 1 0 51244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_553
timestamp 1666464484
transform 1 0 51980 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_557
timestamp 1666464484
transform 1 0 52348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1666464484
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_561
timestamp 1666464484
transform 1 0 52716 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_569
timestamp 1666464484
transform 1 0 53452 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_577
timestamp 1666464484
transform 1 0 54188 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_585
timestamp 1666464484
transform 1 0 54924 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_593
timestamp 1666464484
transform 1 0 55660 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_61_601
timestamp 1666464484
transform 1 0 56396 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_609
timestamp 1666464484
transform 1 0 57132 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_613
timestamp 1666464484
transform 1 0 57500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1666464484
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_61_617
timestamp 1666464484
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_3
timestamp 1666464484
transform 1 0 1380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_11
timestamp 1666464484
transform 1 0 2116 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_19
timestamp 1666464484
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1666464484
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_29
timestamp 1666464484
transform 1 0 3772 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_37
timestamp 1666464484
transform 1 0 4508 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_45
timestamp 1666464484
transform 1 0 5244 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_53
timestamp 1666464484
transform 1 0 5980 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_61
timestamp 1666464484
transform 1 0 6716 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_69
timestamp 1666464484
transform 1 0 7452 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_77
timestamp 1666464484
transform 1 0 8188 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_81
timestamp 1666464484
transform 1 0 8556 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1666464484
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_85
timestamp 1666464484
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_93
timestamp 1666464484
transform 1 0 9660 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_101
timestamp 1666464484
transform 1 0 10396 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_109
timestamp 1666464484
transform 1 0 11132 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_117
timestamp 1666464484
transform 1 0 11868 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_125
timestamp 1666464484
transform 1 0 12604 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_133
timestamp 1666464484
transform 1 0 13340 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_137
timestamp 1666464484
transform 1 0 13708 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1666464484
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_141
timestamp 1666464484
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_149
timestamp 1666464484
transform 1 0 14812 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_157
timestamp 1666464484
transform 1 0 15548 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_165
timestamp 1666464484
transform 1 0 16284 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_173
timestamp 1666464484
transform 1 0 17020 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_181
timestamp 1666464484
transform 1 0 17756 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_189
timestamp 1666464484
transform 1 0 18492 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_193
timestamp 1666464484
transform 1 0 18860 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1666464484
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_197
timestamp 1666464484
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_205
timestamp 1666464484
transform 1 0 19964 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_213
timestamp 1666464484
transform 1 0 20700 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_221
timestamp 1666464484
transform 1 0 21436 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_229
timestamp 1666464484
transform 1 0 22172 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_237
timestamp 1666464484
transform 1 0 22908 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_245
timestamp 1666464484
transform 1 0 23644 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_249
timestamp 1666464484
transform 1 0 24012 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1666464484
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_253
timestamp 1666464484
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_261
timestamp 1666464484
transform 1 0 25116 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_269
timestamp 1666464484
transform 1 0 25852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_277
timestamp 1666464484
transform 1 0 26588 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_285
timestamp 1666464484
transform 1 0 27324 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_293
timestamp 1666464484
transform 1 0 28060 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_301
timestamp 1666464484
transform 1 0 28796 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_305
timestamp 1666464484
transform 1 0 29164 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1666464484
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_309
timestamp 1666464484
transform 1 0 29532 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_317
timestamp 1666464484
transform 1 0 30268 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_325
timestamp 1666464484
transform 1 0 31004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_333
timestamp 1666464484
transform 1 0 31740 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_341
timestamp 1666464484
transform 1 0 32476 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_349
timestamp 1666464484
transform 1 0 33212 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_357
timestamp 1666464484
transform 1 0 33948 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_361
timestamp 1666464484
transform 1 0 34316 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1666464484
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_365
timestamp 1666464484
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_373
timestamp 1666464484
transform 1 0 35420 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_381
timestamp 1666464484
transform 1 0 36156 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_389
timestamp 1666464484
transform 1 0 36892 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_397
timestamp 1666464484
transform 1 0 37628 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_405
timestamp 1666464484
transform 1 0 38364 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_413
timestamp 1666464484
transform 1 0 39100 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_417
timestamp 1666464484
transform 1 0 39468 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1666464484
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_421
timestamp 1666464484
transform 1 0 39836 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_429
timestamp 1666464484
transform 1 0 40572 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_437
timestamp 1666464484
transform 1 0 41308 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_445
timestamp 1666464484
transform 1 0 42044 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_453
timestamp 1666464484
transform 1 0 42780 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_461
timestamp 1666464484
transform 1 0 43516 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_469
timestamp 1666464484
transform 1 0 44252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_473
timestamp 1666464484
transform 1 0 44620 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1666464484
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_477
timestamp 1666464484
transform 1 0 44988 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_485
timestamp 1666464484
transform 1 0 45724 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_493
timestamp 1666464484
transform 1 0 46460 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_501
timestamp 1666464484
transform 1 0 47196 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_509
timestamp 1666464484
transform 1 0 47932 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_517
timestamp 1666464484
transform 1 0 48668 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_525
timestamp 1666464484
transform 1 0 49404 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_529
timestamp 1666464484
transform 1 0 49772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1666464484
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_533
timestamp 1666464484
transform 1 0 50140 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_541
timestamp 1666464484
transform 1 0 50876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_549
timestamp 1666464484
transform 1 0 51612 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_557
timestamp 1666464484
transform 1 0 52348 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_565
timestamp 1666464484
transform 1 0 53084 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_573
timestamp 1666464484
transform 1 0 53820 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_581
timestamp 1666464484
transform 1 0 54556 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_585
timestamp 1666464484
transform 1 0 54924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1666464484
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_589
timestamp 1666464484
transform 1 0 55292 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_597
timestamp 1666464484
transform 1 0 56028 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_605
timestamp 1666464484
transform 1 0 56764 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_62_613
timestamp 1666464484
transform 1 0 57500 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_621
timestamp 1666464484
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_63_3
timestamp 1666464484
transform 1 0 1380 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_11
timestamp 1666464484
transform 1 0 2116 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_19
timestamp 1666464484
transform 1 0 2852 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_27
timestamp 1666464484
transform 1 0 3588 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_35
timestamp 1666464484
transform 1 0 4324 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_43
timestamp 1666464484
transform 1 0 5060 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_51
timestamp 1666464484
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1666464484
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_57
timestamp 1666464484
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_65
timestamp 1666464484
transform 1 0 7084 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_73
timestamp 1666464484
transform 1 0 7820 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_81
timestamp 1666464484
transform 1 0 8556 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_89
timestamp 1666464484
transform 1 0 9292 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_97
timestamp 1666464484
transform 1 0 10028 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_105
timestamp 1666464484
transform 1 0 10764 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_109
timestamp 1666464484
transform 1 0 11132 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1666464484
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_113
timestamp 1666464484
transform 1 0 11500 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_121
timestamp 1666464484
transform 1 0 12236 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_129
timestamp 1666464484
transform 1 0 12972 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_137
timestamp 1666464484
transform 1 0 13708 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_145
timestamp 1666464484
transform 1 0 14444 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_153
timestamp 1666464484
transform 1 0 15180 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_161
timestamp 1666464484
transform 1 0 15916 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_165
timestamp 1666464484
transform 1 0 16284 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1666464484
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_169
timestamp 1666464484
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_177
timestamp 1666464484
transform 1 0 17388 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_185
timestamp 1666464484
transform 1 0 18124 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_193
timestamp 1666464484
transform 1 0 18860 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_201
timestamp 1666464484
transform 1 0 19596 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_209
timestamp 1666464484
transform 1 0 20332 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_217
timestamp 1666464484
transform 1 0 21068 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_221
timestamp 1666464484
transform 1 0 21436 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1666464484
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_225
timestamp 1666464484
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_233
timestamp 1666464484
transform 1 0 22540 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_241
timestamp 1666464484
transform 1 0 23276 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_249
timestamp 1666464484
transform 1 0 24012 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_257
timestamp 1666464484
transform 1 0 24748 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_265
timestamp 1666464484
transform 1 0 25484 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_273
timestamp 1666464484
transform 1 0 26220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_277
timestamp 1666464484
transform 1 0 26588 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1666464484
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_281
timestamp 1666464484
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_289
timestamp 1666464484
transform 1 0 27692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_297
timestamp 1666464484
transform 1 0 28428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_305
timestamp 1666464484
transform 1 0 29164 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_313
timestamp 1666464484
transform 1 0 29900 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_321
timestamp 1666464484
transform 1 0 30636 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_329
timestamp 1666464484
transform 1 0 31372 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_333
timestamp 1666464484
transform 1 0 31740 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1666464484
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_337
timestamp 1666464484
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_345
timestamp 1666464484
transform 1 0 32844 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_353
timestamp 1666464484
transform 1 0 33580 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_361
timestamp 1666464484
transform 1 0 34316 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_369
timestamp 1666464484
transform 1 0 35052 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_377
timestamp 1666464484
transform 1 0 35788 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_385
timestamp 1666464484
transform 1 0 36524 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_389
timestamp 1666464484
transform 1 0 36892 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1666464484
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_393
timestamp 1666464484
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_401
timestamp 1666464484
transform 1 0 37996 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_409
timestamp 1666464484
transform 1 0 38732 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_417
timestamp 1666464484
transform 1 0 39468 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_425
timestamp 1666464484
transform 1 0 40204 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_433
timestamp 1666464484
transform 1 0 40940 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_441
timestamp 1666464484
transform 1 0 41676 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_445
timestamp 1666464484
transform 1 0 42044 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1666464484
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_449
timestamp 1666464484
transform 1 0 42412 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_457
timestamp 1666464484
transform 1 0 43148 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_465
timestamp 1666464484
transform 1 0 43884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_473
timestamp 1666464484
transform 1 0 44620 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_481
timestamp 1666464484
transform 1 0 45356 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_489
timestamp 1666464484
transform 1 0 46092 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_497
timestamp 1666464484
transform 1 0 46828 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_501
timestamp 1666464484
transform 1 0 47196 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1666464484
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_505
timestamp 1666464484
transform 1 0 47564 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_513
timestamp 1666464484
transform 1 0 48300 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_521
timestamp 1666464484
transform 1 0 49036 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_529
timestamp 1666464484
transform 1 0 49772 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_537
timestamp 1666464484
transform 1 0 50508 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_545
timestamp 1666464484
transform 1 0 51244 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_553
timestamp 1666464484
transform 1 0 51980 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_557
timestamp 1666464484
transform 1 0 52348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1666464484
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_561
timestamp 1666464484
transform 1 0 52716 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_569
timestamp 1666464484
transform 1 0 53452 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_577
timestamp 1666464484
transform 1 0 54188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_585
timestamp 1666464484
transform 1 0 54924 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_593
timestamp 1666464484
transform 1 0 55660 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_63_601
timestamp 1666464484
transform 1 0 56396 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_609
timestamp 1666464484
transform 1 0 57132 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_613
timestamp 1666464484
transform 1 0 57500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1666464484
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_63_617
timestamp 1666464484
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_3
timestamp 1666464484
transform 1 0 1380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_11
timestamp 1666464484
transform 1 0 2116 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_19
timestamp 1666464484
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1666464484
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_29
timestamp 1666464484
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_37
timestamp 1666464484
transform 1 0 4508 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_45
timestamp 1666464484
transform 1 0 5244 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_53
timestamp 1666464484
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_61
timestamp 1666464484
transform 1 0 6716 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_69
timestamp 1666464484
transform 1 0 7452 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_77
timestamp 1666464484
transform 1 0 8188 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_81
timestamp 1666464484
transform 1 0 8556 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1666464484
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_85
timestamp 1666464484
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_93
timestamp 1666464484
transform 1 0 9660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_101
timestamp 1666464484
transform 1 0 10396 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_109
timestamp 1666464484
transform 1 0 11132 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_117
timestamp 1666464484
transform 1 0 11868 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_125
timestamp 1666464484
transform 1 0 12604 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_133
timestamp 1666464484
transform 1 0 13340 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_137
timestamp 1666464484
transform 1 0 13708 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1666464484
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_141
timestamp 1666464484
transform 1 0 14076 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_149
timestamp 1666464484
transform 1 0 14812 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_157
timestamp 1666464484
transform 1 0 15548 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_165
timestamp 1666464484
transform 1 0 16284 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_173
timestamp 1666464484
transform 1 0 17020 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_181
timestamp 1666464484
transform 1 0 17756 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_189
timestamp 1666464484
transform 1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_193
timestamp 1666464484
transform 1 0 18860 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1666464484
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_197
timestamp 1666464484
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_205
timestamp 1666464484
transform 1 0 19964 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_213
timestamp 1666464484
transform 1 0 20700 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_221
timestamp 1666464484
transform 1 0 21436 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_229
timestamp 1666464484
transform 1 0 22172 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_237
timestamp 1666464484
transform 1 0 22908 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_245
timestamp 1666464484
transform 1 0 23644 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_249
timestamp 1666464484
transform 1 0 24012 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1666464484
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_253
timestamp 1666464484
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_261
timestamp 1666464484
transform 1 0 25116 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_269
timestamp 1666464484
transform 1 0 25852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_277
timestamp 1666464484
transform 1 0 26588 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_285
timestamp 1666464484
transform 1 0 27324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_293
timestamp 1666464484
transform 1 0 28060 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_301
timestamp 1666464484
transform 1 0 28796 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_305
timestamp 1666464484
transform 1 0 29164 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1666464484
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_309
timestamp 1666464484
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_317
timestamp 1666464484
transform 1 0 30268 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_325
timestamp 1666464484
transform 1 0 31004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_333
timestamp 1666464484
transform 1 0 31740 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_341
timestamp 1666464484
transform 1 0 32476 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_349
timestamp 1666464484
transform 1 0 33212 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_357
timestamp 1666464484
transform 1 0 33948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_361
timestamp 1666464484
transform 1 0 34316 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1666464484
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_365
timestamp 1666464484
transform 1 0 34684 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_373
timestamp 1666464484
transform 1 0 35420 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_381
timestamp 1666464484
transform 1 0 36156 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_389
timestamp 1666464484
transform 1 0 36892 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_397
timestamp 1666464484
transform 1 0 37628 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_405
timestamp 1666464484
transform 1 0 38364 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_413
timestamp 1666464484
transform 1 0 39100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_417
timestamp 1666464484
transform 1 0 39468 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1666464484
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_421
timestamp 1666464484
transform 1 0 39836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_429
timestamp 1666464484
transform 1 0 40572 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_437
timestamp 1666464484
transform 1 0 41308 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_445
timestamp 1666464484
transform 1 0 42044 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_453
timestamp 1666464484
transform 1 0 42780 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_461
timestamp 1666464484
transform 1 0 43516 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_469
timestamp 1666464484
transform 1 0 44252 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_473
timestamp 1666464484
transform 1 0 44620 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1666464484
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_477
timestamp 1666464484
transform 1 0 44988 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_485
timestamp 1666464484
transform 1 0 45724 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_493
timestamp 1666464484
transform 1 0 46460 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_501
timestamp 1666464484
transform 1 0 47196 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_509
timestamp 1666464484
transform 1 0 47932 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_517
timestamp 1666464484
transform 1 0 48668 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_525
timestamp 1666464484
transform 1 0 49404 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_529
timestamp 1666464484
transform 1 0 49772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1666464484
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_533
timestamp 1666464484
transform 1 0 50140 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_541
timestamp 1666464484
transform 1 0 50876 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_549
timestamp 1666464484
transform 1 0 51612 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_557
timestamp 1666464484
transform 1 0 52348 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_565
timestamp 1666464484
transform 1 0 53084 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_573
timestamp 1666464484
transform 1 0 53820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_581
timestamp 1666464484
transform 1 0 54556 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_585
timestamp 1666464484
transform 1 0 54924 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1666464484
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_589
timestamp 1666464484
transform 1 0 55292 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_597
timestamp 1666464484
transform 1 0 56028 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_605
timestamp 1666464484
transform 1 0 56764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_64_613
timestamp 1666464484
transform 1 0 57500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_621
timestamp 1666464484
transform 1 0 58236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_65_3
timestamp 1666464484
transform 1 0 1380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_11
timestamp 1666464484
transform 1 0 2116 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_19
timestamp 1666464484
transform 1 0 2852 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_27
timestamp 1666464484
transform 1 0 3588 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_35
timestamp 1666464484
transform 1 0 4324 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_43
timestamp 1666464484
transform 1 0 5060 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_51
timestamp 1666464484
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1666464484
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_57
timestamp 1666464484
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_65
timestamp 1666464484
transform 1 0 7084 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_73
timestamp 1666464484
transform 1 0 7820 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_81
timestamp 1666464484
transform 1 0 8556 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_89
timestamp 1666464484
transform 1 0 9292 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_97
timestamp 1666464484
transform 1 0 10028 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_105
timestamp 1666464484
transform 1 0 10764 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_109
timestamp 1666464484
transform 1 0 11132 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1666464484
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_113
timestamp 1666464484
transform 1 0 11500 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_121
timestamp 1666464484
transform 1 0 12236 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_129
timestamp 1666464484
transform 1 0 12972 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_137
timestamp 1666464484
transform 1 0 13708 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_145
timestamp 1666464484
transform 1 0 14444 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_153
timestamp 1666464484
transform 1 0 15180 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_161
timestamp 1666464484
transform 1 0 15916 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_165
timestamp 1666464484
transform 1 0 16284 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1666464484
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_169
timestamp 1666464484
transform 1 0 16652 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_177
timestamp 1666464484
transform 1 0 17388 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_185
timestamp 1666464484
transform 1 0 18124 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_193
timestamp 1666464484
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_201
timestamp 1666464484
transform 1 0 19596 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_209
timestamp 1666464484
transform 1 0 20332 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_217
timestamp 1666464484
transform 1 0 21068 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_221
timestamp 1666464484
transform 1 0 21436 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1666464484
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_225
timestamp 1666464484
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_233
timestamp 1666464484
transform 1 0 22540 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_241
timestamp 1666464484
transform 1 0 23276 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_249
timestamp 1666464484
transform 1 0 24012 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_257
timestamp 1666464484
transform 1 0 24748 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_265
timestamp 1666464484
transform 1 0 25484 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_273
timestamp 1666464484
transform 1 0 26220 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_277
timestamp 1666464484
transform 1 0 26588 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1666464484
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_281
timestamp 1666464484
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_289
timestamp 1666464484
transform 1 0 27692 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_297
timestamp 1666464484
transform 1 0 28428 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_305
timestamp 1666464484
transform 1 0 29164 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_313
timestamp 1666464484
transform 1 0 29900 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_321
timestamp 1666464484
transform 1 0 30636 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_329
timestamp 1666464484
transform 1 0 31372 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_333
timestamp 1666464484
transform 1 0 31740 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1666464484
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_337
timestamp 1666464484
transform 1 0 32108 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_345
timestamp 1666464484
transform 1 0 32844 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_353
timestamp 1666464484
transform 1 0 33580 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_361
timestamp 1666464484
transform 1 0 34316 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_369
timestamp 1666464484
transform 1 0 35052 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_377
timestamp 1666464484
transform 1 0 35788 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_385
timestamp 1666464484
transform 1 0 36524 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_389
timestamp 1666464484
transform 1 0 36892 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1666464484
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_393
timestamp 1666464484
transform 1 0 37260 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_401
timestamp 1666464484
transform 1 0 37996 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_409
timestamp 1666464484
transform 1 0 38732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_417
timestamp 1666464484
transform 1 0 39468 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_425
timestamp 1666464484
transform 1 0 40204 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_433
timestamp 1666464484
transform 1 0 40940 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_441
timestamp 1666464484
transform 1 0 41676 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_445
timestamp 1666464484
transform 1 0 42044 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1666464484
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_449
timestamp 1666464484
transform 1 0 42412 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_457
timestamp 1666464484
transform 1 0 43148 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_465
timestamp 1666464484
transform 1 0 43884 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_473
timestamp 1666464484
transform 1 0 44620 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_481
timestamp 1666464484
transform 1 0 45356 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_489
timestamp 1666464484
transform 1 0 46092 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_497
timestamp 1666464484
transform 1 0 46828 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_501
timestamp 1666464484
transform 1 0 47196 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1666464484
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_505
timestamp 1666464484
transform 1 0 47564 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_513
timestamp 1666464484
transform 1 0 48300 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_521
timestamp 1666464484
transform 1 0 49036 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_529
timestamp 1666464484
transform 1 0 49772 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_537
timestamp 1666464484
transform 1 0 50508 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_545
timestamp 1666464484
transform 1 0 51244 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_553
timestamp 1666464484
transform 1 0 51980 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_557
timestamp 1666464484
transform 1 0 52348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1666464484
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_561
timestamp 1666464484
transform 1 0 52716 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_569
timestamp 1666464484
transform 1 0 53452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_577
timestamp 1666464484
transform 1 0 54188 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_585
timestamp 1666464484
transform 1 0 54924 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_593
timestamp 1666464484
transform 1 0 55660 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_65_601
timestamp 1666464484
transform 1 0 56396 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_609
timestamp 1666464484
transform 1 0 57132 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_613
timestamp 1666464484
transform 1 0 57500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1666464484
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_617
timestamp 1666464484
transform 1 0 57868 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_3
timestamp 1666464484
transform 1 0 1380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_11
timestamp 1666464484
transform 1 0 2116 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_19
timestamp 1666464484
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1666464484
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_29
timestamp 1666464484
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_37
timestamp 1666464484
transform 1 0 4508 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_45
timestamp 1666464484
transform 1 0 5244 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_53
timestamp 1666464484
transform 1 0 5980 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_61
timestamp 1666464484
transform 1 0 6716 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_69
timestamp 1666464484
transform 1 0 7452 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_77
timestamp 1666464484
transform 1 0 8188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_81
timestamp 1666464484
transform 1 0 8556 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1666464484
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_85
timestamp 1666464484
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_93
timestamp 1666464484
transform 1 0 9660 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_101
timestamp 1666464484
transform 1 0 10396 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_109
timestamp 1666464484
transform 1 0 11132 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_117
timestamp 1666464484
transform 1 0 11868 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_125
timestamp 1666464484
transform 1 0 12604 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_133
timestamp 1666464484
transform 1 0 13340 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_137
timestamp 1666464484
transform 1 0 13708 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1666464484
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_141
timestamp 1666464484
transform 1 0 14076 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_149
timestamp 1666464484
transform 1 0 14812 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_157
timestamp 1666464484
transform 1 0 15548 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_165
timestamp 1666464484
transform 1 0 16284 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_173
timestamp 1666464484
transform 1 0 17020 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_181
timestamp 1666464484
transform 1 0 17756 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_189
timestamp 1666464484
transform 1 0 18492 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_193
timestamp 1666464484
transform 1 0 18860 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1666464484
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_197
timestamp 1666464484
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_205
timestamp 1666464484
transform 1 0 19964 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_213
timestamp 1666464484
transform 1 0 20700 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_221
timestamp 1666464484
transform 1 0 21436 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_229
timestamp 1666464484
transform 1 0 22172 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_237
timestamp 1666464484
transform 1 0 22908 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_245
timestamp 1666464484
transform 1 0 23644 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_249
timestamp 1666464484
transform 1 0 24012 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1666464484
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_253
timestamp 1666464484
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_261
timestamp 1666464484
transform 1 0 25116 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_269
timestamp 1666464484
transform 1 0 25852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_277
timestamp 1666464484
transform 1 0 26588 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_285
timestamp 1666464484
transform 1 0 27324 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_293
timestamp 1666464484
transform 1 0 28060 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_301
timestamp 1666464484
transform 1 0 28796 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_305
timestamp 1666464484
transform 1 0 29164 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1666464484
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_309
timestamp 1666464484
transform 1 0 29532 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_317
timestamp 1666464484
transform 1 0 30268 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_325
timestamp 1666464484
transform 1 0 31004 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_333
timestamp 1666464484
transform 1 0 31740 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_341
timestamp 1666464484
transform 1 0 32476 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_349
timestamp 1666464484
transform 1 0 33212 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_357
timestamp 1666464484
transform 1 0 33948 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_361
timestamp 1666464484
transform 1 0 34316 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1666464484
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_365
timestamp 1666464484
transform 1 0 34684 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_373
timestamp 1666464484
transform 1 0 35420 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_381
timestamp 1666464484
transform 1 0 36156 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_389
timestamp 1666464484
transform 1 0 36892 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_397
timestamp 1666464484
transform 1 0 37628 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_405
timestamp 1666464484
transform 1 0 38364 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_413
timestamp 1666464484
transform 1 0 39100 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_417
timestamp 1666464484
transform 1 0 39468 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1666464484
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_421
timestamp 1666464484
transform 1 0 39836 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_429
timestamp 1666464484
transform 1 0 40572 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_437
timestamp 1666464484
transform 1 0 41308 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_445
timestamp 1666464484
transform 1 0 42044 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_453
timestamp 1666464484
transform 1 0 42780 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_461
timestamp 1666464484
transform 1 0 43516 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_469
timestamp 1666464484
transform 1 0 44252 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_473
timestamp 1666464484
transform 1 0 44620 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1666464484
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_477
timestamp 1666464484
transform 1 0 44988 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_485
timestamp 1666464484
transform 1 0 45724 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_493
timestamp 1666464484
transform 1 0 46460 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_501
timestamp 1666464484
transform 1 0 47196 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_509
timestamp 1666464484
transform 1 0 47932 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_517
timestamp 1666464484
transform 1 0 48668 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_525
timestamp 1666464484
transform 1 0 49404 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_529
timestamp 1666464484
transform 1 0 49772 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1666464484
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_533
timestamp 1666464484
transform 1 0 50140 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_541
timestamp 1666464484
transform 1 0 50876 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_549
timestamp 1666464484
transform 1 0 51612 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_557
timestamp 1666464484
transform 1 0 52348 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_565
timestamp 1666464484
transform 1 0 53084 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_573
timestamp 1666464484
transform 1 0 53820 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_581
timestamp 1666464484
transform 1 0 54556 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_585
timestamp 1666464484
transform 1 0 54924 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1666464484
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_589
timestamp 1666464484
transform 1 0 55292 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_597
timestamp 1666464484
transform 1 0 56028 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_605
timestamp 1666464484
transform 1 0 56764 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_66_613
timestamp 1666464484
transform 1 0 57500 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_621
timestamp 1666464484
transform 1 0 58236 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_67_3
timestamp 1666464484
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_11
timestamp 1666464484
transform 1 0 2116 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_19
timestamp 1666464484
transform 1 0 2852 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_27
timestamp 1666464484
transform 1 0 3588 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_35
timestamp 1666464484
transform 1 0 4324 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_43
timestamp 1666464484
transform 1 0 5060 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_51
timestamp 1666464484
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1666464484
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_57
timestamp 1666464484
transform 1 0 6348 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_65
timestamp 1666464484
transform 1 0 7084 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_73
timestamp 1666464484
transform 1 0 7820 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_81
timestamp 1666464484
transform 1 0 8556 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_89
timestamp 1666464484
transform 1 0 9292 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_97
timestamp 1666464484
transform 1 0 10028 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_105
timestamp 1666464484
transform 1 0 10764 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_109
timestamp 1666464484
transform 1 0 11132 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1666464484
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_113
timestamp 1666464484
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_121
timestamp 1666464484
transform 1 0 12236 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_129
timestamp 1666464484
transform 1 0 12972 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_137
timestamp 1666464484
transform 1 0 13708 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_145
timestamp 1666464484
transform 1 0 14444 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_153
timestamp 1666464484
transform 1 0 15180 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_161
timestamp 1666464484
transform 1 0 15916 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_165
timestamp 1666464484
transform 1 0 16284 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1666464484
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_169
timestamp 1666464484
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_177
timestamp 1666464484
transform 1 0 17388 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_185
timestamp 1666464484
transform 1 0 18124 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_193
timestamp 1666464484
transform 1 0 18860 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_201
timestamp 1666464484
transform 1 0 19596 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_209
timestamp 1666464484
transform 1 0 20332 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_217
timestamp 1666464484
transform 1 0 21068 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_221
timestamp 1666464484
transform 1 0 21436 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1666464484
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_225
timestamp 1666464484
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_233
timestamp 1666464484
transform 1 0 22540 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_241
timestamp 1666464484
transform 1 0 23276 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_249
timestamp 1666464484
transform 1 0 24012 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_257
timestamp 1666464484
transform 1 0 24748 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_265
timestamp 1666464484
transform 1 0 25484 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_273
timestamp 1666464484
transform 1 0 26220 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_277
timestamp 1666464484
transform 1 0 26588 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1666464484
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_281
timestamp 1666464484
transform 1 0 26956 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_289
timestamp 1666464484
transform 1 0 27692 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_297
timestamp 1666464484
transform 1 0 28428 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_305
timestamp 1666464484
transform 1 0 29164 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_313
timestamp 1666464484
transform 1 0 29900 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_321
timestamp 1666464484
transform 1 0 30636 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_329
timestamp 1666464484
transform 1 0 31372 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_333
timestamp 1666464484
transform 1 0 31740 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1666464484
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_337
timestamp 1666464484
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_345
timestamp 1666464484
transform 1 0 32844 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_353
timestamp 1666464484
transform 1 0 33580 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_361
timestamp 1666464484
transform 1 0 34316 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_369
timestamp 1666464484
transform 1 0 35052 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_377
timestamp 1666464484
transform 1 0 35788 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_385
timestamp 1666464484
transform 1 0 36524 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_389
timestamp 1666464484
transform 1 0 36892 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1666464484
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_393
timestamp 1666464484
transform 1 0 37260 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_401
timestamp 1666464484
transform 1 0 37996 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_409
timestamp 1666464484
transform 1 0 38732 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_417
timestamp 1666464484
transform 1 0 39468 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_425
timestamp 1666464484
transform 1 0 40204 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_433
timestamp 1666464484
transform 1 0 40940 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_441
timestamp 1666464484
transform 1 0 41676 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_445
timestamp 1666464484
transform 1 0 42044 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1666464484
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_449
timestamp 1666464484
transform 1 0 42412 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_457
timestamp 1666464484
transform 1 0 43148 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_465
timestamp 1666464484
transform 1 0 43884 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_473
timestamp 1666464484
transform 1 0 44620 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_481
timestamp 1666464484
transform 1 0 45356 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_489
timestamp 1666464484
transform 1 0 46092 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_497
timestamp 1666464484
transform 1 0 46828 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_501
timestamp 1666464484
transform 1 0 47196 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1666464484
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_505
timestamp 1666464484
transform 1 0 47564 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_513
timestamp 1666464484
transform 1 0 48300 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_521
timestamp 1666464484
transform 1 0 49036 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_529
timestamp 1666464484
transform 1 0 49772 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_537
timestamp 1666464484
transform 1 0 50508 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_545
timestamp 1666464484
transform 1 0 51244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_553
timestamp 1666464484
transform 1 0 51980 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_557
timestamp 1666464484
transform 1 0 52348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1666464484
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_561
timestamp 1666464484
transform 1 0 52716 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_569
timestamp 1666464484
transform 1 0 53452 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_577
timestamp 1666464484
transform 1 0 54188 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_585
timestamp 1666464484
transform 1 0 54924 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_593
timestamp 1666464484
transform 1 0 55660 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_67_601
timestamp 1666464484
transform 1 0 56396 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_609
timestamp 1666464484
transform 1 0 57132 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_613
timestamp 1666464484
transform 1 0 57500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1666464484
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_617
timestamp 1666464484
transform 1 0 57868 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_3
timestamp 1666464484
transform 1 0 1380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_11
timestamp 1666464484
transform 1 0 2116 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_19
timestamp 1666464484
transform 1 0 2852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1666464484
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_29
timestamp 1666464484
transform 1 0 3772 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_37
timestamp 1666464484
transform 1 0 4508 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_45
timestamp 1666464484
transform 1 0 5244 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_53
timestamp 1666464484
transform 1 0 5980 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_61
timestamp 1666464484
transform 1 0 6716 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_69
timestamp 1666464484
transform 1 0 7452 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_77
timestamp 1666464484
transform 1 0 8188 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_81
timestamp 1666464484
transform 1 0 8556 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1666464484
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_85
timestamp 1666464484
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_93
timestamp 1666464484
transform 1 0 9660 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_101
timestamp 1666464484
transform 1 0 10396 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_109
timestamp 1666464484
transform 1 0 11132 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_117
timestamp 1666464484
transform 1 0 11868 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_125
timestamp 1666464484
transform 1 0 12604 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_133
timestamp 1666464484
transform 1 0 13340 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_137
timestamp 1666464484
transform 1 0 13708 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1666464484
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_141
timestamp 1666464484
transform 1 0 14076 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_149
timestamp 1666464484
transform 1 0 14812 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_157
timestamp 1666464484
transform 1 0 15548 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_165
timestamp 1666464484
transform 1 0 16284 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_173
timestamp 1666464484
transform 1 0 17020 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_181
timestamp 1666464484
transform 1 0 17756 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_189
timestamp 1666464484
transform 1 0 18492 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_193
timestamp 1666464484
transform 1 0 18860 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1666464484
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_197
timestamp 1666464484
transform 1 0 19228 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_205
timestamp 1666464484
transform 1 0 19964 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_213
timestamp 1666464484
transform 1 0 20700 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_221
timestamp 1666464484
transform 1 0 21436 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_229
timestamp 1666464484
transform 1 0 22172 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_237
timestamp 1666464484
transform 1 0 22908 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_245
timestamp 1666464484
transform 1 0 23644 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_249
timestamp 1666464484
transform 1 0 24012 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1666464484
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_253
timestamp 1666464484
transform 1 0 24380 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_261
timestamp 1666464484
transform 1 0 25116 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_269
timestamp 1666464484
transform 1 0 25852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_277
timestamp 1666464484
transform 1 0 26588 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_285
timestamp 1666464484
transform 1 0 27324 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_293
timestamp 1666464484
transform 1 0 28060 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_301
timestamp 1666464484
transform 1 0 28796 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_305
timestamp 1666464484
transform 1 0 29164 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1666464484
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_309
timestamp 1666464484
transform 1 0 29532 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_317
timestamp 1666464484
transform 1 0 30268 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_325
timestamp 1666464484
transform 1 0 31004 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_333
timestamp 1666464484
transform 1 0 31740 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_341
timestamp 1666464484
transform 1 0 32476 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_349
timestamp 1666464484
transform 1 0 33212 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_357
timestamp 1666464484
transform 1 0 33948 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_361
timestamp 1666464484
transform 1 0 34316 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1666464484
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_365
timestamp 1666464484
transform 1 0 34684 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_373
timestamp 1666464484
transform 1 0 35420 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_381
timestamp 1666464484
transform 1 0 36156 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_389
timestamp 1666464484
transform 1 0 36892 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_397
timestamp 1666464484
transform 1 0 37628 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_405
timestamp 1666464484
transform 1 0 38364 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_413
timestamp 1666464484
transform 1 0 39100 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_417
timestamp 1666464484
transform 1 0 39468 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1666464484
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_421
timestamp 1666464484
transform 1 0 39836 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_429
timestamp 1666464484
transform 1 0 40572 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_437
timestamp 1666464484
transform 1 0 41308 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_445
timestamp 1666464484
transform 1 0 42044 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_453
timestamp 1666464484
transform 1 0 42780 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_461
timestamp 1666464484
transform 1 0 43516 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_469
timestamp 1666464484
transform 1 0 44252 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_473
timestamp 1666464484
transform 1 0 44620 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1666464484
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_477
timestamp 1666464484
transform 1 0 44988 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_485
timestamp 1666464484
transform 1 0 45724 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_493
timestamp 1666464484
transform 1 0 46460 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_501
timestamp 1666464484
transform 1 0 47196 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_509
timestamp 1666464484
transform 1 0 47932 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_517
timestamp 1666464484
transform 1 0 48668 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_525
timestamp 1666464484
transform 1 0 49404 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_529
timestamp 1666464484
transform 1 0 49772 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1666464484
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_533
timestamp 1666464484
transform 1 0 50140 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_541
timestamp 1666464484
transform 1 0 50876 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_549
timestamp 1666464484
transform 1 0 51612 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_557
timestamp 1666464484
transform 1 0 52348 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_565
timestamp 1666464484
transform 1 0 53084 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_573
timestamp 1666464484
transform 1 0 53820 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_581
timestamp 1666464484
transform 1 0 54556 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_585
timestamp 1666464484
transform 1 0 54924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1666464484
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_68_589
timestamp 1666464484
transform 1 0 55292 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_597
timestamp 1666464484
transform 1 0 56028 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_605
timestamp 1666464484
transform 1 0 56764 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_68_613
timestamp 1666464484
transform 1 0 57500 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_68_621
timestamp 1666464484
transform 1 0 58236 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_69_3
timestamp 1666464484
transform 1 0 1380 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_11
timestamp 1666464484
transform 1 0 2116 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_19
timestamp 1666464484
transform 1 0 2852 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_27
timestamp 1666464484
transform 1 0 3588 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_35
timestamp 1666464484
transform 1 0 4324 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_43
timestamp 1666464484
transform 1 0 5060 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_51
timestamp 1666464484
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1666464484
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_57
timestamp 1666464484
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_65
timestamp 1666464484
transform 1 0 7084 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_73
timestamp 1666464484
transform 1 0 7820 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_81
timestamp 1666464484
transform 1 0 8556 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_89
timestamp 1666464484
transform 1 0 9292 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_97
timestamp 1666464484
transform 1 0 10028 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_105
timestamp 1666464484
transform 1 0 10764 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_109
timestamp 1666464484
transform 1 0 11132 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1666464484
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_113
timestamp 1666464484
transform 1 0 11500 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_121
timestamp 1666464484
transform 1 0 12236 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_129
timestamp 1666464484
transform 1 0 12972 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_137
timestamp 1666464484
transform 1 0 13708 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_145
timestamp 1666464484
transform 1 0 14444 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_153
timestamp 1666464484
transform 1 0 15180 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_161
timestamp 1666464484
transform 1 0 15916 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_165
timestamp 1666464484
transform 1 0 16284 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1666464484
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_169
timestamp 1666464484
transform 1 0 16652 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_177
timestamp 1666464484
transform 1 0 17388 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_185
timestamp 1666464484
transform 1 0 18124 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_193
timestamp 1666464484
transform 1 0 18860 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_201
timestamp 1666464484
transform 1 0 19596 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_209
timestamp 1666464484
transform 1 0 20332 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_217
timestamp 1666464484
transform 1 0 21068 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_221
timestamp 1666464484
transform 1 0 21436 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1666464484
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_225
timestamp 1666464484
transform 1 0 21804 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_233
timestamp 1666464484
transform 1 0 22540 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_241
timestamp 1666464484
transform 1 0 23276 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_249
timestamp 1666464484
transform 1 0 24012 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_257
timestamp 1666464484
transform 1 0 24748 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_265
timestamp 1666464484
transform 1 0 25484 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_273
timestamp 1666464484
transform 1 0 26220 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_277
timestamp 1666464484
transform 1 0 26588 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1666464484
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_281
timestamp 1666464484
transform 1 0 26956 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_289
timestamp 1666464484
transform 1 0 27692 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_297
timestamp 1666464484
transform 1 0 28428 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_305
timestamp 1666464484
transform 1 0 29164 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_313
timestamp 1666464484
transform 1 0 29900 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_321
timestamp 1666464484
transform 1 0 30636 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_329
timestamp 1666464484
transform 1 0 31372 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_333
timestamp 1666464484
transform 1 0 31740 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1666464484
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_337
timestamp 1666464484
transform 1 0 32108 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_345
timestamp 1666464484
transform 1 0 32844 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_353
timestamp 1666464484
transform 1 0 33580 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_361
timestamp 1666464484
transform 1 0 34316 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_369
timestamp 1666464484
transform 1 0 35052 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_377
timestamp 1666464484
transform 1 0 35788 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_385
timestamp 1666464484
transform 1 0 36524 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_389
timestamp 1666464484
transform 1 0 36892 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1666464484
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_393
timestamp 1666464484
transform 1 0 37260 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_401
timestamp 1666464484
transform 1 0 37996 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_409
timestamp 1666464484
transform 1 0 38732 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_417
timestamp 1666464484
transform 1 0 39468 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_425
timestamp 1666464484
transform 1 0 40204 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_433
timestamp 1666464484
transform 1 0 40940 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_441
timestamp 1666464484
transform 1 0 41676 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_445
timestamp 1666464484
transform 1 0 42044 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1666464484
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_449
timestamp 1666464484
transform 1 0 42412 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_457
timestamp 1666464484
transform 1 0 43148 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_465
timestamp 1666464484
transform 1 0 43884 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_473
timestamp 1666464484
transform 1 0 44620 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_481
timestamp 1666464484
transform 1 0 45356 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_489
timestamp 1666464484
transform 1 0 46092 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_497
timestamp 1666464484
transform 1 0 46828 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_501
timestamp 1666464484
transform 1 0 47196 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1666464484
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_505
timestamp 1666464484
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_513
timestamp 1666464484
transform 1 0 48300 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_521
timestamp 1666464484
transform 1 0 49036 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_529
timestamp 1666464484
transform 1 0 49772 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_537
timestamp 1666464484
transform 1 0 50508 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_545
timestamp 1666464484
transform 1 0 51244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_553
timestamp 1666464484
transform 1 0 51980 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_557
timestamp 1666464484
transform 1 0 52348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1666464484
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_561
timestamp 1666464484
transform 1 0 52716 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_569
timestamp 1666464484
transform 1 0 53452 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_577
timestamp 1666464484
transform 1 0 54188 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_585
timestamp 1666464484
transform 1 0 54924 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_593
timestamp 1666464484
transform 1 0 55660 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_69_601
timestamp 1666464484
transform 1 0 56396 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_69_609
timestamp 1666464484
transform 1 0 57132 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_613
timestamp 1666464484
transform 1 0 57500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1666464484
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_69_617
timestamp 1666464484
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_3
timestamp 1666464484
transform 1 0 1380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_11
timestamp 1666464484
transform 1 0 2116 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_19
timestamp 1666464484
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1666464484
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_29
timestamp 1666464484
transform 1 0 3772 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_37
timestamp 1666464484
transform 1 0 4508 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_45
timestamp 1666464484
transform 1 0 5244 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_53
timestamp 1666464484
transform 1 0 5980 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_61
timestamp 1666464484
transform 1 0 6716 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_69
timestamp 1666464484
transform 1 0 7452 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_77
timestamp 1666464484
transform 1 0 8188 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_81
timestamp 1666464484
transform 1 0 8556 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1666464484
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_85
timestamp 1666464484
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_93
timestamp 1666464484
transform 1 0 9660 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_101
timestamp 1666464484
transform 1 0 10396 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_109
timestamp 1666464484
transform 1 0 11132 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_117
timestamp 1666464484
transform 1 0 11868 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_125
timestamp 1666464484
transform 1 0 12604 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_133
timestamp 1666464484
transform 1 0 13340 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_137
timestamp 1666464484
transform 1 0 13708 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1666464484
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_141
timestamp 1666464484
transform 1 0 14076 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_149
timestamp 1666464484
transform 1 0 14812 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_157
timestamp 1666464484
transform 1 0 15548 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_165
timestamp 1666464484
transform 1 0 16284 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_173
timestamp 1666464484
transform 1 0 17020 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_181
timestamp 1666464484
transform 1 0 17756 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_189
timestamp 1666464484
transform 1 0 18492 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_193
timestamp 1666464484
transform 1 0 18860 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1666464484
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_197
timestamp 1666464484
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_205
timestamp 1666464484
transform 1 0 19964 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_213
timestamp 1666464484
transform 1 0 20700 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_221
timestamp 1666464484
transform 1 0 21436 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_229
timestamp 1666464484
transform 1 0 22172 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_237
timestamp 1666464484
transform 1 0 22908 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_245
timestamp 1666464484
transform 1 0 23644 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_249
timestamp 1666464484
transform 1 0 24012 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1666464484
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_253
timestamp 1666464484
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_261
timestamp 1666464484
transform 1 0 25116 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_269
timestamp 1666464484
transform 1 0 25852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_277
timestamp 1666464484
transform 1 0 26588 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_285
timestamp 1666464484
transform 1 0 27324 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_293
timestamp 1666464484
transform 1 0 28060 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_301
timestamp 1666464484
transform 1 0 28796 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_305
timestamp 1666464484
transform 1 0 29164 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1666464484
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_309
timestamp 1666464484
transform 1 0 29532 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_317
timestamp 1666464484
transform 1 0 30268 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_325
timestamp 1666464484
transform 1 0 31004 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_333
timestamp 1666464484
transform 1 0 31740 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_341
timestamp 1666464484
transform 1 0 32476 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_349
timestamp 1666464484
transform 1 0 33212 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_357
timestamp 1666464484
transform 1 0 33948 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_361
timestamp 1666464484
transform 1 0 34316 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1666464484
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_365
timestamp 1666464484
transform 1 0 34684 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_373
timestamp 1666464484
transform 1 0 35420 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_381
timestamp 1666464484
transform 1 0 36156 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_389
timestamp 1666464484
transform 1 0 36892 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_397
timestamp 1666464484
transform 1 0 37628 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_405
timestamp 1666464484
transform 1 0 38364 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_413
timestamp 1666464484
transform 1 0 39100 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_417
timestamp 1666464484
transform 1 0 39468 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1666464484
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_421
timestamp 1666464484
transform 1 0 39836 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_429
timestamp 1666464484
transform 1 0 40572 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_437
timestamp 1666464484
transform 1 0 41308 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_445
timestamp 1666464484
transform 1 0 42044 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_453
timestamp 1666464484
transform 1 0 42780 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_461
timestamp 1666464484
transform 1 0 43516 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_469
timestamp 1666464484
transform 1 0 44252 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_473
timestamp 1666464484
transform 1 0 44620 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1666464484
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_477
timestamp 1666464484
transform 1 0 44988 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_485
timestamp 1666464484
transform 1 0 45724 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_493
timestamp 1666464484
transform 1 0 46460 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_501
timestamp 1666464484
transform 1 0 47196 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_509
timestamp 1666464484
transform 1 0 47932 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_517
timestamp 1666464484
transform 1 0 48668 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_525
timestamp 1666464484
transform 1 0 49404 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_529
timestamp 1666464484
transform 1 0 49772 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1666464484
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_533
timestamp 1666464484
transform 1 0 50140 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_541
timestamp 1666464484
transform 1 0 50876 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_549
timestamp 1666464484
transform 1 0 51612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_557
timestamp 1666464484
transform 1 0 52348 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_565
timestamp 1666464484
transform 1 0 53084 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_573
timestamp 1666464484
transform 1 0 53820 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_581
timestamp 1666464484
transform 1 0 54556 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_585
timestamp 1666464484
transform 1 0 54924 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1666464484
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_589
timestamp 1666464484
transform 1 0 55292 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_597
timestamp 1666464484
transform 1 0 56028 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_605
timestamp 1666464484
transform 1 0 56764 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_613
timestamp 1666464484
transform 1 0 57500 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_621
timestamp 1666464484
transform 1 0 58236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_71_3
timestamp 1666464484
transform 1 0 1380 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_11
timestamp 1666464484
transform 1 0 2116 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_19
timestamp 1666464484
transform 1 0 2852 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_27
timestamp 1666464484
transform 1 0 3588 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_35
timestamp 1666464484
transform 1 0 4324 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_43
timestamp 1666464484
transform 1 0 5060 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_51
timestamp 1666464484
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1666464484
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_57
timestamp 1666464484
transform 1 0 6348 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_65
timestamp 1666464484
transform 1 0 7084 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_73
timestamp 1666464484
transform 1 0 7820 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_81
timestamp 1666464484
transform 1 0 8556 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_89
timestamp 1666464484
transform 1 0 9292 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_97
timestamp 1666464484
transform 1 0 10028 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_105
timestamp 1666464484
transform 1 0 10764 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_109
timestamp 1666464484
transform 1 0 11132 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1666464484
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_113
timestamp 1666464484
transform 1 0 11500 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_121
timestamp 1666464484
transform 1 0 12236 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_129
timestamp 1666464484
transform 1 0 12972 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_137
timestamp 1666464484
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_145
timestamp 1666464484
transform 1 0 14444 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_153
timestamp 1666464484
transform 1 0 15180 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_161
timestamp 1666464484
transform 1 0 15916 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_165
timestamp 1666464484
transform 1 0 16284 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1666464484
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_169
timestamp 1666464484
transform 1 0 16652 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_177
timestamp 1666464484
transform 1 0 17388 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_185
timestamp 1666464484
transform 1 0 18124 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_193
timestamp 1666464484
transform 1 0 18860 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_201
timestamp 1666464484
transform 1 0 19596 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_209
timestamp 1666464484
transform 1 0 20332 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_217
timestamp 1666464484
transform 1 0 21068 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_221
timestamp 1666464484
transform 1 0 21436 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1666464484
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_225
timestamp 1666464484
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_233
timestamp 1666464484
transform 1 0 22540 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_241
timestamp 1666464484
transform 1 0 23276 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_249
timestamp 1666464484
transform 1 0 24012 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_257
timestamp 1666464484
transform 1 0 24748 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_265
timestamp 1666464484
transform 1 0 25484 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_273
timestamp 1666464484
transform 1 0 26220 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_277
timestamp 1666464484
transform 1 0 26588 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1666464484
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_281
timestamp 1666464484
transform 1 0 26956 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_289
timestamp 1666464484
transform 1 0 27692 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_297
timestamp 1666464484
transform 1 0 28428 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_305
timestamp 1666464484
transform 1 0 29164 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_313
timestamp 1666464484
transform 1 0 29900 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_321
timestamp 1666464484
transform 1 0 30636 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_329
timestamp 1666464484
transform 1 0 31372 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_333
timestamp 1666464484
transform 1 0 31740 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1666464484
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_337
timestamp 1666464484
transform 1 0 32108 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_345
timestamp 1666464484
transform 1 0 32844 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_353
timestamp 1666464484
transform 1 0 33580 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_361
timestamp 1666464484
transform 1 0 34316 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_369
timestamp 1666464484
transform 1 0 35052 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_377
timestamp 1666464484
transform 1 0 35788 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_385
timestamp 1666464484
transform 1 0 36524 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_389
timestamp 1666464484
transform 1 0 36892 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1666464484
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_393
timestamp 1666464484
transform 1 0 37260 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_401
timestamp 1666464484
transform 1 0 37996 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_409
timestamp 1666464484
transform 1 0 38732 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_417
timestamp 1666464484
transform 1 0 39468 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_425
timestamp 1666464484
transform 1 0 40204 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_433
timestamp 1666464484
transform 1 0 40940 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_441
timestamp 1666464484
transform 1 0 41676 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_445
timestamp 1666464484
transform 1 0 42044 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1666464484
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_449
timestamp 1666464484
transform 1 0 42412 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_457
timestamp 1666464484
transform 1 0 43148 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_465
timestamp 1666464484
transform 1 0 43884 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_473
timestamp 1666464484
transform 1 0 44620 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_481
timestamp 1666464484
transform 1 0 45356 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_489
timestamp 1666464484
transform 1 0 46092 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_497
timestamp 1666464484
transform 1 0 46828 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_501
timestamp 1666464484
transform 1 0 47196 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1666464484
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_505
timestamp 1666464484
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_513
timestamp 1666464484
transform 1 0 48300 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_521
timestamp 1666464484
transform 1 0 49036 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_529
timestamp 1666464484
transform 1 0 49772 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_537
timestamp 1666464484
transform 1 0 50508 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_545
timestamp 1666464484
transform 1 0 51244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_553
timestamp 1666464484
transform 1 0 51980 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_557
timestamp 1666464484
transform 1 0 52348 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1666464484
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_561
timestamp 1666464484
transform 1 0 52716 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_569
timestamp 1666464484
transform 1 0 53452 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_577
timestamp 1666464484
transform 1 0 54188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_585
timestamp 1666464484
transform 1 0 54924 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_593
timestamp 1666464484
transform 1 0 55660 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_71_601
timestamp 1666464484
transform 1 0 56396 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_609
timestamp 1666464484
transform 1 0 57132 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_613
timestamp 1666464484
transform 1 0 57500 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1666464484
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_71_617
timestamp 1666464484
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_3
timestamp 1666464484
transform 1 0 1380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_11
timestamp 1666464484
transform 1 0 2116 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_19
timestamp 1666464484
transform 1 0 2852 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1666464484
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_29
timestamp 1666464484
transform 1 0 3772 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_37
timestamp 1666464484
transform 1 0 4508 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_45
timestamp 1666464484
transform 1 0 5244 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_53
timestamp 1666464484
transform 1 0 5980 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_61
timestamp 1666464484
transform 1 0 6716 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_69
timestamp 1666464484
transform 1 0 7452 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_77
timestamp 1666464484
transform 1 0 8188 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_81
timestamp 1666464484
transform 1 0 8556 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1666464484
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_85
timestamp 1666464484
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_93
timestamp 1666464484
transform 1 0 9660 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_101
timestamp 1666464484
transform 1 0 10396 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_109
timestamp 1666464484
transform 1 0 11132 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_117
timestamp 1666464484
transform 1 0 11868 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_125
timestamp 1666464484
transform 1 0 12604 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_133
timestamp 1666464484
transform 1 0 13340 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_137
timestamp 1666464484
transform 1 0 13708 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1666464484
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_141
timestamp 1666464484
transform 1 0 14076 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_149
timestamp 1666464484
transform 1 0 14812 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_157
timestamp 1666464484
transform 1 0 15548 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_165
timestamp 1666464484
transform 1 0 16284 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_173
timestamp 1666464484
transform 1 0 17020 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_181
timestamp 1666464484
transform 1 0 17756 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_189
timestamp 1666464484
transform 1 0 18492 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_193
timestamp 1666464484
transform 1 0 18860 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1666464484
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_197
timestamp 1666464484
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_205
timestamp 1666464484
transform 1 0 19964 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_213
timestamp 1666464484
transform 1 0 20700 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_221
timestamp 1666464484
transform 1 0 21436 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_229
timestamp 1666464484
transform 1 0 22172 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_237
timestamp 1666464484
transform 1 0 22908 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_245
timestamp 1666464484
transform 1 0 23644 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_249
timestamp 1666464484
transform 1 0 24012 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1666464484
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_253
timestamp 1666464484
transform 1 0 24380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_261
timestamp 1666464484
transform 1 0 25116 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_269
timestamp 1666464484
transform 1 0 25852 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_277
timestamp 1666464484
transform 1 0 26588 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_285
timestamp 1666464484
transform 1 0 27324 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_293
timestamp 1666464484
transform 1 0 28060 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_301
timestamp 1666464484
transform 1 0 28796 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_305
timestamp 1666464484
transform 1 0 29164 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1666464484
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_309
timestamp 1666464484
transform 1 0 29532 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_317
timestamp 1666464484
transform 1 0 30268 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_325
timestamp 1666464484
transform 1 0 31004 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_333
timestamp 1666464484
transform 1 0 31740 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_341
timestamp 1666464484
transform 1 0 32476 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_349
timestamp 1666464484
transform 1 0 33212 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_357
timestamp 1666464484
transform 1 0 33948 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_361
timestamp 1666464484
transform 1 0 34316 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1666464484
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_365
timestamp 1666464484
transform 1 0 34684 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_373
timestamp 1666464484
transform 1 0 35420 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_381
timestamp 1666464484
transform 1 0 36156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_389
timestamp 1666464484
transform 1 0 36892 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_397
timestamp 1666464484
transform 1 0 37628 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_405
timestamp 1666464484
transform 1 0 38364 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_413
timestamp 1666464484
transform 1 0 39100 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_417
timestamp 1666464484
transform 1 0 39468 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1666464484
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_421
timestamp 1666464484
transform 1 0 39836 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_429
timestamp 1666464484
transform 1 0 40572 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_437
timestamp 1666464484
transform 1 0 41308 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_445
timestamp 1666464484
transform 1 0 42044 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_453
timestamp 1666464484
transform 1 0 42780 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_461
timestamp 1666464484
transform 1 0 43516 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_469
timestamp 1666464484
transform 1 0 44252 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_473
timestamp 1666464484
transform 1 0 44620 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1666464484
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_477
timestamp 1666464484
transform 1 0 44988 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_485
timestamp 1666464484
transform 1 0 45724 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_493
timestamp 1666464484
transform 1 0 46460 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_501
timestamp 1666464484
transform 1 0 47196 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_509
timestamp 1666464484
transform 1 0 47932 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_517
timestamp 1666464484
transform 1 0 48668 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_525
timestamp 1666464484
transform 1 0 49404 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_529
timestamp 1666464484
transform 1 0 49772 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1666464484
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_533
timestamp 1666464484
transform 1 0 50140 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_541
timestamp 1666464484
transform 1 0 50876 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_549
timestamp 1666464484
transform 1 0 51612 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_557
timestamp 1666464484
transform 1 0 52348 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_565
timestamp 1666464484
transform 1 0 53084 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_573
timestamp 1666464484
transform 1 0 53820 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_581
timestamp 1666464484
transform 1 0 54556 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_585
timestamp 1666464484
transform 1 0 54924 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1666464484
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_589
timestamp 1666464484
transform 1 0 55292 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_597
timestamp 1666464484
transform 1 0 56028 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_605
timestamp 1666464484
transform 1 0 56764 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_72_613
timestamp 1666464484
transform 1 0 57500 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_72_621
timestamp 1666464484
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_73_3
timestamp 1666464484
transform 1 0 1380 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_11
timestamp 1666464484
transform 1 0 2116 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_19
timestamp 1666464484
transform 1 0 2852 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_27
timestamp 1666464484
transform 1 0 3588 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_35
timestamp 1666464484
transform 1 0 4324 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_43
timestamp 1666464484
transform 1 0 5060 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_51
timestamp 1666464484
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1666464484
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_57
timestamp 1666464484
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_65
timestamp 1666464484
transform 1 0 7084 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_73
timestamp 1666464484
transform 1 0 7820 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_81
timestamp 1666464484
transform 1 0 8556 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_89
timestamp 1666464484
transform 1 0 9292 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_97
timestamp 1666464484
transform 1 0 10028 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_105
timestamp 1666464484
transform 1 0 10764 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_109
timestamp 1666464484
transform 1 0 11132 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1666464484
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_113
timestamp 1666464484
transform 1 0 11500 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_121
timestamp 1666464484
transform 1 0 12236 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_129
timestamp 1666464484
transform 1 0 12972 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_137
timestamp 1666464484
transform 1 0 13708 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_145
timestamp 1666464484
transform 1 0 14444 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_153
timestamp 1666464484
transform 1 0 15180 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_161
timestamp 1666464484
transform 1 0 15916 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_165
timestamp 1666464484
transform 1 0 16284 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1666464484
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_169
timestamp 1666464484
transform 1 0 16652 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_177
timestamp 1666464484
transform 1 0 17388 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_185
timestamp 1666464484
transform 1 0 18124 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_193
timestamp 1666464484
transform 1 0 18860 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_201
timestamp 1666464484
transform 1 0 19596 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_209
timestamp 1666464484
transform 1 0 20332 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_217
timestamp 1666464484
transform 1 0 21068 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_221
timestamp 1666464484
transform 1 0 21436 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1666464484
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_225
timestamp 1666464484
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_233
timestamp 1666464484
transform 1 0 22540 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_241
timestamp 1666464484
transform 1 0 23276 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_249
timestamp 1666464484
transform 1 0 24012 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_257
timestamp 1666464484
transform 1 0 24748 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_265
timestamp 1666464484
transform 1 0 25484 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_273
timestamp 1666464484
transform 1 0 26220 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_277
timestamp 1666464484
transform 1 0 26588 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1666464484
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_281
timestamp 1666464484
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_289
timestamp 1666464484
transform 1 0 27692 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_297
timestamp 1666464484
transform 1 0 28428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_305
timestamp 1666464484
transform 1 0 29164 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_313
timestamp 1666464484
transform 1 0 29900 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_321
timestamp 1666464484
transform 1 0 30636 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_329
timestamp 1666464484
transform 1 0 31372 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_333
timestamp 1666464484
transform 1 0 31740 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1666464484
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_337
timestamp 1666464484
transform 1 0 32108 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_345
timestamp 1666464484
transform 1 0 32844 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_353
timestamp 1666464484
transform 1 0 33580 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_361
timestamp 1666464484
transform 1 0 34316 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_369
timestamp 1666464484
transform 1 0 35052 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_377
timestamp 1666464484
transform 1 0 35788 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_385
timestamp 1666464484
transform 1 0 36524 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_389
timestamp 1666464484
transform 1 0 36892 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1666464484
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_393
timestamp 1666464484
transform 1 0 37260 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_401
timestamp 1666464484
transform 1 0 37996 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_409
timestamp 1666464484
transform 1 0 38732 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_417
timestamp 1666464484
transform 1 0 39468 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_425
timestamp 1666464484
transform 1 0 40204 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_433
timestamp 1666464484
transform 1 0 40940 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_441
timestamp 1666464484
transform 1 0 41676 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_445
timestamp 1666464484
transform 1 0 42044 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1666464484
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_449
timestamp 1666464484
transform 1 0 42412 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_457
timestamp 1666464484
transform 1 0 43148 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_465
timestamp 1666464484
transform 1 0 43884 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_473
timestamp 1666464484
transform 1 0 44620 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_481
timestamp 1666464484
transform 1 0 45356 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_489
timestamp 1666464484
transform 1 0 46092 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_497
timestamp 1666464484
transform 1 0 46828 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_501
timestamp 1666464484
transform 1 0 47196 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1666464484
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_505
timestamp 1666464484
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_513
timestamp 1666464484
transform 1 0 48300 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_521
timestamp 1666464484
transform 1 0 49036 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_529
timestamp 1666464484
transform 1 0 49772 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_537
timestamp 1666464484
transform 1 0 50508 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_545
timestamp 1666464484
transform 1 0 51244 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_553
timestamp 1666464484
transform 1 0 51980 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_557
timestamp 1666464484
transform 1 0 52348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1666464484
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_561
timestamp 1666464484
transform 1 0 52716 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_569
timestamp 1666464484
transform 1 0 53452 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_577
timestamp 1666464484
transform 1 0 54188 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_585
timestamp 1666464484
transform 1 0 54924 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_593
timestamp 1666464484
transform 1 0 55660 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_601
timestamp 1666464484
transform 1 0 56396 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_73_609
timestamp 1666464484
transform 1 0 57132 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_613
timestamp 1666464484
transform 1 0 57500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1666464484
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_73_617
timestamp 1666464484
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_3
timestamp 1666464484
transform 1 0 1380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_11
timestamp 1666464484
transform 1 0 2116 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_19
timestamp 1666464484
transform 1 0 2852 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1666464484
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_29
timestamp 1666464484
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_37
timestamp 1666464484
transform 1 0 4508 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_45
timestamp 1666464484
transform 1 0 5244 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_53
timestamp 1666464484
transform 1 0 5980 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_61
timestamp 1666464484
transform 1 0 6716 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_69
timestamp 1666464484
transform 1 0 7452 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_77
timestamp 1666464484
transform 1 0 8188 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_81
timestamp 1666464484
transform 1 0 8556 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1666464484
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_85
timestamp 1666464484
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_93
timestamp 1666464484
transform 1 0 9660 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_101
timestamp 1666464484
transform 1 0 10396 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_109
timestamp 1666464484
transform 1 0 11132 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_117
timestamp 1666464484
transform 1 0 11868 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_125
timestamp 1666464484
transform 1 0 12604 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_133
timestamp 1666464484
transform 1 0 13340 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_137
timestamp 1666464484
transform 1 0 13708 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1666464484
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_141
timestamp 1666464484
transform 1 0 14076 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_149
timestamp 1666464484
transform 1 0 14812 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_157
timestamp 1666464484
transform 1 0 15548 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_165
timestamp 1666464484
transform 1 0 16284 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_173
timestamp 1666464484
transform 1 0 17020 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_181
timestamp 1666464484
transform 1 0 17756 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_189
timestamp 1666464484
transform 1 0 18492 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_193
timestamp 1666464484
transform 1 0 18860 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1666464484
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_197
timestamp 1666464484
transform 1 0 19228 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_205
timestamp 1666464484
transform 1 0 19964 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_213
timestamp 1666464484
transform 1 0 20700 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_221
timestamp 1666464484
transform 1 0 21436 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_229
timestamp 1666464484
transform 1 0 22172 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_237
timestamp 1666464484
transform 1 0 22908 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_245
timestamp 1666464484
transform 1 0 23644 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_249
timestamp 1666464484
transform 1 0 24012 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1666464484
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_253
timestamp 1666464484
transform 1 0 24380 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_261
timestamp 1666464484
transform 1 0 25116 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_269
timestamp 1666464484
transform 1 0 25852 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_277
timestamp 1666464484
transform 1 0 26588 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_285
timestamp 1666464484
transform 1 0 27324 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_293
timestamp 1666464484
transform 1 0 28060 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_301
timestamp 1666464484
transform 1 0 28796 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_305
timestamp 1666464484
transform 1 0 29164 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1666464484
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_309
timestamp 1666464484
transform 1 0 29532 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_317
timestamp 1666464484
transform 1 0 30268 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_325
timestamp 1666464484
transform 1 0 31004 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_333
timestamp 1666464484
transform 1 0 31740 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_341
timestamp 1666464484
transform 1 0 32476 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_349
timestamp 1666464484
transform 1 0 33212 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_357
timestamp 1666464484
transform 1 0 33948 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_361
timestamp 1666464484
transform 1 0 34316 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1666464484
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_365
timestamp 1666464484
transform 1 0 34684 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_373
timestamp 1666464484
transform 1 0 35420 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_381
timestamp 1666464484
transform 1 0 36156 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_389
timestamp 1666464484
transform 1 0 36892 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_397
timestamp 1666464484
transform 1 0 37628 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_405
timestamp 1666464484
transform 1 0 38364 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_413
timestamp 1666464484
transform 1 0 39100 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_417
timestamp 1666464484
transform 1 0 39468 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1666464484
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_421
timestamp 1666464484
transform 1 0 39836 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_429
timestamp 1666464484
transform 1 0 40572 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_437
timestamp 1666464484
transform 1 0 41308 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_445
timestamp 1666464484
transform 1 0 42044 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_453
timestamp 1666464484
transform 1 0 42780 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_461
timestamp 1666464484
transform 1 0 43516 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_469
timestamp 1666464484
transform 1 0 44252 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_473
timestamp 1666464484
transform 1 0 44620 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1666464484
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_477
timestamp 1666464484
transform 1 0 44988 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_485
timestamp 1666464484
transform 1 0 45724 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_493
timestamp 1666464484
transform 1 0 46460 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_501
timestamp 1666464484
transform 1 0 47196 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_509
timestamp 1666464484
transform 1 0 47932 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_517
timestamp 1666464484
transform 1 0 48668 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_525
timestamp 1666464484
transform 1 0 49404 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_529
timestamp 1666464484
transform 1 0 49772 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1666464484
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_533
timestamp 1666464484
transform 1 0 50140 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_541
timestamp 1666464484
transform 1 0 50876 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_549
timestamp 1666464484
transform 1 0 51612 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_557
timestamp 1666464484
transform 1 0 52348 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_565
timestamp 1666464484
transform 1 0 53084 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_573
timestamp 1666464484
transform 1 0 53820 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_581
timestamp 1666464484
transform 1 0 54556 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_585
timestamp 1666464484
transform 1 0 54924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1666464484
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_74_589
timestamp 1666464484
transform 1 0 55292 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_597
timestamp 1666464484
transform 1 0 56028 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_605
timestamp 1666464484
transform 1 0 56764 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_74_613
timestamp 1666464484
transform 1 0 57500 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_74_621
timestamp 1666464484
transform 1 0 58236 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_75_3
timestamp 1666464484
transform 1 0 1380 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_11
timestamp 1666464484
transform 1 0 2116 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_19
timestamp 1666464484
transform 1 0 2852 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_27
timestamp 1666464484
transform 1 0 3588 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_35
timestamp 1666464484
transform 1 0 4324 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_43
timestamp 1666464484
transform 1 0 5060 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_51
timestamp 1666464484
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1666464484
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_57
timestamp 1666464484
transform 1 0 6348 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_65
timestamp 1666464484
transform 1 0 7084 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_73
timestamp 1666464484
transform 1 0 7820 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_81
timestamp 1666464484
transform 1 0 8556 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_89
timestamp 1666464484
transform 1 0 9292 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_97
timestamp 1666464484
transform 1 0 10028 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_105
timestamp 1666464484
transform 1 0 10764 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_109
timestamp 1666464484
transform 1 0 11132 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1666464484
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_113
timestamp 1666464484
transform 1 0 11500 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_121
timestamp 1666464484
transform 1 0 12236 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_129
timestamp 1666464484
transform 1 0 12972 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_137
timestamp 1666464484
transform 1 0 13708 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_145
timestamp 1666464484
transform 1 0 14444 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_153
timestamp 1666464484
transform 1 0 15180 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_161
timestamp 1666464484
transform 1 0 15916 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_165
timestamp 1666464484
transform 1 0 16284 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1666464484
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_169
timestamp 1666464484
transform 1 0 16652 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_177
timestamp 1666464484
transform 1 0 17388 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_185
timestamp 1666464484
transform 1 0 18124 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_193
timestamp 1666464484
transform 1 0 18860 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_201
timestamp 1666464484
transform 1 0 19596 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_209
timestamp 1666464484
transform 1 0 20332 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_217
timestamp 1666464484
transform 1 0 21068 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_221
timestamp 1666464484
transform 1 0 21436 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1666464484
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_225
timestamp 1666464484
transform 1 0 21804 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_233
timestamp 1666464484
transform 1 0 22540 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_241
timestamp 1666464484
transform 1 0 23276 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_249
timestamp 1666464484
transform 1 0 24012 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_257
timestamp 1666464484
transform 1 0 24748 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_265
timestamp 1666464484
transform 1 0 25484 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_273
timestamp 1666464484
transform 1 0 26220 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_277
timestamp 1666464484
transform 1 0 26588 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1666464484
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_281
timestamp 1666464484
transform 1 0 26956 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_289
timestamp 1666464484
transform 1 0 27692 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_297
timestamp 1666464484
transform 1 0 28428 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_305
timestamp 1666464484
transform 1 0 29164 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_313
timestamp 1666464484
transform 1 0 29900 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_321
timestamp 1666464484
transform 1 0 30636 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_329
timestamp 1666464484
transform 1 0 31372 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_333
timestamp 1666464484
transform 1 0 31740 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1666464484
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_337
timestamp 1666464484
transform 1 0 32108 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_345
timestamp 1666464484
transform 1 0 32844 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_353
timestamp 1666464484
transform 1 0 33580 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_361
timestamp 1666464484
transform 1 0 34316 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_369
timestamp 1666464484
transform 1 0 35052 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_377
timestamp 1666464484
transform 1 0 35788 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_385
timestamp 1666464484
transform 1 0 36524 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_389
timestamp 1666464484
transform 1 0 36892 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1666464484
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_393
timestamp 1666464484
transform 1 0 37260 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_401
timestamp 1666464484
transform 1 0 37996 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_409
timestamp 1666464484
transform 1 0 38732 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_417
timestamp 1666464484
transform 1 0 39468 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_425
timestamp 1666464484
transform 1 0 40204 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_433
timestamp 1666464484
transform 1 0 40940 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_441
timestamp 1666464484
transform 1 0 41676 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_445
timestamp 1666464484
transform 1 0 42044 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1666464484
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_449
timestamp 1666464484
transform 1 0 42412 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_457
timestamp 1666464484
transform 1 0 43148 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_465
timestamp 1666464484
transform 1 0 43884 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_473
timestamp 1666464484
transform 1 0 44620 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_481
timestamp 1666464484
transform 1 0 45356 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_489
timestamp 1666464484
transform 1 0 46092 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_497
timestamp 1666464484
transform 1 0 46828 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_501
timestamp 1666464484
transform 1 0 47196 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1666464484
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_505
timestamp 1666464484
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_513
timestamp 1666464484
transform 1 0 48300 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_521
timestamp 1666464484
transform 1 0 49036 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_529
timestamp 1666464484
transform 1 0 49772 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_537
timestamp 1666464484
transform 1 0 50508 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_545
timestamp 1666464484
transform 1 0 51244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_553
timestamp 1666464484
transform 1 0 51980 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_557
timestamp 1666464484
transform 1 0 52348 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1666464484
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_561
timestamp 1666464484
transform 1 0 52716 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_569
timestamp 1666464484
transform 1 0 53452 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_577
timestamp 1666464484
transform 1 0 54188 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_585
timestamp 1666464484
transform 1 0 54924 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_593
timestamp 1666464484
transform 1 0 55660 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_75_601
timestamp 1666464484
transform 1 0 56396 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_609
timestamp 1666464484
transform 1 0 57132 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_613
timestamp 1666464484
transform 1 0 57500 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1666464484
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_617
timestamp 1666464484
transform 1 0 57868 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_3
timestamp 1666464484
transform 1 0 1380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_11
timestamp 1666464484
transform 1 0 2116 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_19
timestamp 1666464484
transform 1 0 2852 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1666464484
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_29
timestamp 1666464484
transform 1 0 3772 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_37
timestamp 1666464484
transform 1 0 4508 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_45
timestamp 1666464484
transform 1 0 5244 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_53
timestamp 1666464484
transform 1 0 5980 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_61
timestamp 1666464484
transform 1 0 6716 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_69
timestamp 1666464484
transform 1 0 7452 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_77
timestamp 1666464484
transform 1 0 8188 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_81
timestamp 1666464484
transform 1 0 8556 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1666464484
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_85
timestamp 1666464484
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_93
timestamp 1666464484
transform 1 0 9660 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_101
timestamp 1666464484
transform 1 0 10396 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_109
timestamp 1666464484
transform 1 0 11132 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_117
timestamp 1666464484
transform 1 0 11868 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_125
timestamp 1666464484
transform 1 0 12604 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_133
timestamp 1666464484
transform 1 0 13340 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_137
timestamp 1666464484
transform 1 0 13708 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1666464484
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_141
timestamp 1666464484
transform 1 0 14076 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_149
timestamp 1666464484
transform 1 0 14812 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_157
timestamp 1666464484
transform 1 0 15548 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_165
timestamp 1666464484
transform 1 0 16284 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_173
timestamp 1666464484
transform 1 0 17020 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_181
timestamp 1666464484
transform 1 0 17756 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_189
timestamp 1666464484
transform 1 0 18492 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_193
timestamp 1666464484
transform 1 0 18860 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1666464484
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_197
timestamp 1666464484
transform 1 0 19228 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_205
timestamp 1666464484
transform 1 0 19964 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_213
timestamp 1666464484
transform 1 0 20700 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_221
timestamp 1666464484
transform 1 0 21436 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_229
timestamp 1666464484
transform 1 0 22172 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_237
timestamp 1666464484
transform 1 0 22908 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_245
timestamp 1666464484
transform 1 0 23644 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_249
timestamp 1666464484
transform 1 0 24012 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1666464484
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_253
timestamp 1666464484
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_261
timestamp 1666464484
transform 1 0 25116 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_269
timestamp 1666464484
transform 1 0 25852 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_277
timestamp 1666464484
transform 1 0 26588 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_285
timestamp 1666464484
transform 1 0 27324 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_293
timestamp 1666464484
transform 1 0 28060 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_301
timestamp 1666464484
transform 1 0 28796 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_305
timestamp 1666464484
transform 1 0 29164 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1666464484
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_309
timestamp 1666464484
transform 1 0 29532 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_317
timestamp 1666464484
transform 1 0 30268 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_325
timestamp 1666464484
transform 1 0 31004 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_333
timestamp 1666464484
transform 1 0 31740 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_341
timestamp 1666464484
transform 1 0 32476 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_349
timestamp 1666464484
transform 1 0 33212 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_357
timestamp 1666464484
transform 1 0 33948 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_361
timestamp 1666464484
transform 1 0 34316 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1666464484
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_365
timestamp 1666464484
transform 1 0 34684 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_373
timestamp 1666464484
transform 1 0 35420 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_381
timestamp 1666464484
transform 1 0 36156 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_389
timestamp 1666464484
transform 1 0 36892 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_397
timestamp 1666464484
transform 1 0 37628 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_405
timestamp 1666464484
transform 1 0 38364 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_413
timestamp 1666464484
transform 1 0 39100 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_417
timestamp 1666464484
transform 1 0 39468 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1666464484
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_421
timestamp 1666464484
transform 1 0 39836 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_429
timestamp 1666464484
transform 1 0 40572 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_437
timestamp 1666464484
transform 1 0 41308 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_445
timestamp 1666464484
transform 1 0 42044 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_453
timestamp 1666464484
transform 1 0 42780 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_461
timestamp 1666464484
transform 1 0 43516 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_469
timestamp 1666464484
transform 1 0 44252 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_473
timestamp 1666464484
transform 1 0 44620 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1666464484
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_477
timestamp 1666464484
transform 1 0 44988 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_485
timestamp 1666464484
transform 1 0 45724 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_493
timestamp 1666464484
transform 1 0 46460 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_501
timestamp 1666464484
transform 1 0 47196 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_509
timestamp 1666464484
transform 1 0 47932 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_517
timestamp 1666464484
transform 1 0 48668 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_525
timestamp 1666464484
transform 1 0 49404 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_529
timestamp 1666464484
transform 1 0 49772 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1666464484
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_533
timestamp 1666464484
transform 1 0 50140 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_541
timestamp 1666464484
transform 1 0 50876 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_549
timestamp 1666464484
transform 1 0 51612 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_557
timestamp 1666464484
transform 1 0 52348 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_565
timestamp 1666464484
transform 1 0 53084 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_573
timestamp 1666464484
transform 1 0 53820 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_581
timestamp 1666464484
transform 1 0 54556 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_585
timestamp 1666464484
transform 1 0 54924 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1666464484
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_76_589
timestamp 1666464484
transform 1 0 55292 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_597
timestamp 1666464484
transform 1 0 56028 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_605
timestamp 1666464484
transform 1 0 56764 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_76_613
timestamp 1666464484
transform 1 0 57500 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_76_621
timestamp 1666464484
transform 1 0 58236 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_77_3
timestamp 1666464484
transform 1 0 1380 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_11
timestamp 1666464484
transform 1 0 2116 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_19
timestamp 1666464484
transform 1 0 2852 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_27
timestamp 1666464484
transform 1 0 3588 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_35
timestamp 1666464484
transform 1 0 4324 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_43
timestamp 1666464484
transform 1 0 5060 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_51
timestamp 1666464484
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1666464484
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_57
timestamp 1666464484
transform 1 0 6348 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_65
timestamp 1666464484
transform 1 0 7084 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_73
timestamp 1666464484
transform 1 0 7820 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_81
timestamp 1666464484
transform 1 0 8556 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_89
timestamp 1666464484
transform 1 0 9292 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_97
timestamp 1666464484
transform 1 0 10028 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_105
timestamp 1666464484
transform 1 0 10764 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_109
timestamp 1666464484
transform 1 0 11132 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1666464484
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_113
timestamp 1666464484
transform 1 0 11500 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_121
timestamp 1666464484
transform 1 0 12236 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_129
timestamp 1666464484
transform 1 0 12972 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_137
timestamp 1666464484
transform 1 0 13708 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_145
timestamp 1666464484
transform 1 0 14444 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_153
timestamp 1666464484
transform 1 0 15180 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_161
timestamp 1666464484
transform 1 0 15916 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_165
timestamp 1666464484
transform 1 0 16284 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1666464484
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_169
timestamp 1666464484
transform 1 0 16652 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_177
timestamp 1666464484
transform 1 0 17388 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_185
timestamp 1666464484
transform 1 0 18124 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_193
timestamp 1666464484
transform 1 0 18860 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_201
timestamp 1666464484
transform 1 0 19596 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_209
timestamp 1666464484
transform 1 0 20332 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_217
timestamp 1666464484
transform 1 0 21068 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_221
timestamp 1666464484
transform 1 0 21436 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1666464484
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_225
timestamp 1666464484
transform 1 0 21804 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_233
timestamp 1666464484
transform 1 0 22540 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_241
timestamp 1666464484
transform 1 0 23276 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_249
timestamp 1666464484
transform 1 0 24012 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_257
timestamp 1666464484
transform 1 0 24748 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_265
timestamp 1666464484
transform 1 0 25484 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_273
timestamp 1666464484
transform 1 0 26220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_277
timestamp 1666464484
transform 1 0 26588 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1666464484
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_281
timestamp 1666464484
transform 1 0 26956 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_289
timestamp 1666464484
transform 1 0 27692 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_297
timestamp 1666464484
transform 1 0 28428 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_305
timestamp 1666464484
transform 1 0 29164 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_313
timestamp 1666464484
transform 1 0 29900 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_321
timestamp 1666464484
transform 1 0 30636 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_329
timestamp 1666464484
transform 1 0 31372 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_333
timestamp 1666464484
transform 1 0 31740 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1666464484
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_337
timestamp 1666464484
transform 1 0 32108 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_345
timestamp 1666464484
transform 1 0 32844 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_353
timestamp 1666464484
transform 1 0 33580 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_361
timestamp 1666464484
transform 1 0 34316 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_369
timestamp 1666464484
transform 1 0 35052 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_377
timestamp 1666464484
transform 1 0 35788 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_385
timestamp 1666464484
transform 1 0 36524 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_389
timestamp 1666464484
transform 1 0 36892 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1666464484
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_393
timestamp 1666464484
transform 1 0 37260 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_401
timestamp 1666464484
transform 1 0 37996 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_409
timestamp 1666464484
transform 1 0 38732 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_417
timestamp 1666464484
transform 1 0 39468 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_425
timestamp 1666464484
transform 1 0 40204 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_433
timestamp 1666464484
transform 1 0 40940 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_441
timestamp 1666464484
transform 1 0 41676 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_445
timestamp 1666464484
transform 1 0 42044 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1666464484
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_449
timestamp 1666464484
transform 1 0 42412 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_457
timestamp 1666464484
transform 1 0 43148 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_465
timestamp 1666464484
transform 1 0 43884 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_473
timestamp 1666464484
transform 1 0 44620 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_481
timestamp 1666464484
transform 1 0 45356 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_489
timestamp 1666464484
transform 1 0 46092 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_497
timestamp 1666464484
transform 1 0 46828 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_501
timestamp 1666464484
transform 1 0 47196 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1666464484
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_505
timestamp 1666464484
transform 1 0 47564 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_513
timestamp 1666464484
transform 1 0 48300 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_521
timestamp 1666464484
transform 1 0 49036 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_529
timestamp 1666464484
transform 1 0 49772 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_537
timestamp 1666464484
transform 1 0 50508 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_545
timestamp 1666464484
transform 1 0 51244 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_553
timestamp 1666464484
transform 1 0 51980 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_557
timestamp 1666464484
transform 1 0 52348 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1666464484
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_561
timestamp 1666464484
transform 1 0 52716 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_569
timestamp 1666464484
transform 1 0 53452 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_577
timestamp 1666464484
transform 1 0 54188 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_585
timestamp 1666464484
transform 1 0 54924 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_593
timestamp 1666464484
transform 1 0 55660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_77_601
timestamp 1666464484
transform 1 0 56396 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_77_609
timestamp 1666464484
transform 1 0 57132 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_613
timestamp 1666464484
transform 1 0 57500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1666464484
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_77_617
timestamp 1666464484
transform 1 0 57868 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_3
timestamp 1666464484
transform 1 0 1380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_11
timestamp 1666464484
transform 1 0 2116 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_19
timestamp 1666464484
transform 1 0 2852 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1666464484
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_29
timestamp 1666464484
transform 1 0 3772 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_37
timestamp 1666464484
transform 1 0 4508 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_45
timestamp 1666464484
transform 1 0 5244 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_53
timestamp 1666464484
transform 1 0 5980 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_61
timestamp 1666464484
transform 1 0 6716 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_69
timestamp 1666464484
transform 1 0 7452 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_77
timestamp 1666464484
transform 1 0 8188 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_81
timestamp 1666464484
transform 1 0 8556 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1666464484
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_85
timestamp 1666464484
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_93
timestamp 1666464484
transform 1 0 9660 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_101
timestamp 1666464484
transform 1 0 10396 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_109
timestamp 1666464484
transform 1 0 11132 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_117
timestamp 1666464484
transform 1 0 11868 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_125
timestamp 1666464484
transform 1 0 12604 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_133
timestamp 1666464484
transform 1 0 13340 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_137
timestamp 1666464484
transform 1 0 13708 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1666464484
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_141
timestamp 1666464484
transform 1 0 14076 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_149
timestamp 1666464484
transform 1 0 14812 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_157
timestamp 1666464484
transform 1 0 15548 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_165
timestamp 1666464484
transform 1 0 16284 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_173
timestamp 1666464484
transform 1 0 17020 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_181
timestamp 1666464484
transform 1 0 17756 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_189
timestamp 1666464484
transform 1 0 18492 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_193
timestamp 1666464484
transform 1 0 18860 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1666464484
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_197
timestamp 1666464484
transform 1 0 19228 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_205
timestamp 1666464484
transform 1 0 19964 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_213
timestamp 1666464484
transform 1 0 20700 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_221
timestamp 1666464484
transform 1 0 21436 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_229
timestamp 1666464484
transform 1 0 22172 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_237
timestamp 1666464484
transform 1 0 22908 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_245
timestamp 1666464484
transform 1 0 23644 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_249
timestamp 1666464484
transform 1 0 24012 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1666464484
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_253
timestamp 1666464484
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_261
timestamp 1666464484
transform 1 0 25116 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_269
timestamp 1666464484
transform 1 0 25852 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_277
timestamp 1666464484
transform 1 0 26588 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_285
timestamp 1666464484
transform 1 0 27324 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_293
timestamp 1666464484
transform 1 0 28060 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_301
timestamp 1666464484
transform 1 0 28796 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_305
timestamp 1666464484
transform 1 0 29164 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1666464484
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_309
timestamp 1666464484
transform 1 0 29532 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_317
timestamp 1666464484
transform 1 0 30268 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_325
timestamp 1666464484
transform 1 0 31004 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_333
timestamp 1666464484
transform 1 0 31740 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_341
timestamp 1666464484
transform 1 0 32476 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_349
timestamp 1666464484
transform 1 0 33212 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_357
timestamp 1666464484
transform 1 0 33948 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_361
timestamp 1666464484
transform 1 0 34316 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1666464484
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_365
timestamp 1666464484
transform 1 0 34684 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_373
timestamp 1666464484
transform 1 0 35420 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_381
timestamp 1666464484
transform 1 0 36156 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_389
timestamp 1666464484
transform 1 0 36892 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_397
timestamp 1666464484
transform 1 0 37628 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_405
timestamp 1666464484
transform 1 0 38364 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_413
timestamp 1666464484
transform 1 0 39100 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_417
timestamp 1666464484
transform 1 0 39468 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1666464484
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_421
timestamp 1666464484
transform 1 0 39836 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_429
timestamp 1666464484
transform 1 0 40572 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_437
timestamp 1666464484
transform 1 0 41308 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_445
timestamp 1666464484
transform 1 0 42044 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_453
timestamp 1666464484
transform 1 0 42780 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_461
timestamp 1666464484
transform 1 0 43516 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_469
timestamp 1666464484
transform 1 0 44252 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_473
timestamp 1666464484
transform 1 0 44620 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1666464484
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_477
timestamp 1666464484
transform 1 0 44988 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_485
timestamp 1666464484
transform 1 0 45724 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_493
timestamp 1666464484
transform 1 0 46460 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_501
timestamp 1666464484
transform 1 0 47196 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_509
timestamp 1666464484
transform 1 0 47932 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_517
timestamp 1666464484
transform 1 0 48668 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_525
timestamp 1666464484
transform 1 0 49404 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_529
timestamp 1666464484
transform 1 0 49772 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1666464484
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_533
timestamp 1666464484
transform 1 0 50140 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_541
timestamp 1666464484
transform 1 0 50876 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_549
timestamp 1666464484
transform 1 0 51612 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_557
timestamp 1666464484
transform 1 0 52348 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_565
timestamp 1666464484
transform 1 0 53084 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_573
timestamp 1666464484
transform 1 0 53820 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_581
timestamp 1666464484
transform 1 0 54556 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_585
timestamp 1666464484
transform 1 0 54924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1666464484
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_78_589
timestamp 1666464484
transform 1 0 55292 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_597
timestamp 1666464484
transform 1 0 56028 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_605
timestamp 1666464484
transform 1 0 56764 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_78_613
timestamp 1666464484
transform 1 0 57500 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_78_621
timestamp 1666464484
transform 1 0 58236 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_79_3
timestamp 1666464484
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_11
timestamp 1666464484
transform 1 0 2116 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_19
timestamp 1666464484
transform 1 0 2852 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_27
timestamp 1666464484
transform 1 0 3588 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_35
timestamp 1666464484
transform 1 0 4324 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_43
timestamp 1666464484
transform 1 0 5060 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_51
timestamp 1666464484
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1666464484
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_57
timestamp 1666464484
transform 1 0 6348 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_65
timestamp 1666464484
transform 1 0 7084 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_73
timestamp 1666464484
transform 1 0 7820 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_81
timestamp 1666464484
transform 1 0 8556 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_89
timestamp 1666464484
transform 1 0 9292 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_97
timestamp 1666464484
transform 1 0 10028 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_105
timestamp 1666464484
transform 1 0 10764 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_109
timestamp 1666464484
transform 1 0 11132 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1666464484
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_113
timestamp 1666464484
transform 1 0 11500 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_121
timestamp 1666464484
transform 1 0 12236 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_129
timestamp 1666464484
transform 1 0 12972 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_137
timestamp 1666464484
transform 1 0 13708 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_145
timestamp 1666464484
transform 1 0 14444 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_153
timestamp 1666464484
transform 1 0 15180 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_161
timestamp 1666464484
transform 1 0 15916 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_165
timestamp 1666464484
transform 1 0 16284 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1666464484
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_169
timestamp 1666464484
transform 1 0 16652 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_177
timestamp 1666464484
transform 1 0 17388 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_185
timestamp 1666464484
transform 1 0 18124 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_193
timestamp 1666464484
transform 1 0 18860 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_201
timestamp 1666464484
transform 1 0 19596 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_209
timestamp 1666464484
transform 1 0 20332 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_217
timestamp 1666464484
transform 1 0 21068 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_221
timestamp 1666464484
transform 1 0 21436 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1666464484
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_225
timestamp 1666464484
transform 1 0 21804 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_233
timestamp 1666464484
transform 1 0 22540 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_241
timestamp 1666464484
transform 1 0 23276 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_249
timestamp 1666464484
transform 1 0 24012 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_257
timestamp 1666464484
transform 1 0 24748 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_265
timestamp 1666464484
transform 1 0 25484 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_273
timestamp 1666464484
transform 1 0 26220 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_277
timestamp 1666464484
transform 1 0 26588 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1666464484
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_281
timestamp 1666464484
transform 1 0 26956 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_289
timestamp 1666464484
transform 1 0 27692 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_297
timestamp 1666464484
transform 1 0 28428 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_305
timestamp 1666464484
transform 1 0 29164 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_313
timestamp 1666464484
transform 1 0 29900 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_321
timestamp 1666464484
transform 1 0 30636 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_329
timestamp 1666464484
transform 1 0 31372 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_333
timestamp 1666464484
transform 1 0 31740 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1666464484
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_337
timestamp 1666464484
transform 1 0 32108 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_345
timestamp 1666464484
transform 1 0 32844 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_353
timestamp 1666464484
transform 1 0 33580 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_361
timestamp 1666464484
transform 1 0 34316 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_369
timestamp 1666464484
transform 1 0 35052 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_377
timestamp 1666464484
transform 1 0 35788 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_385
timestamp 1666464484
transform 1 0 36524 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_389
timestamp 1666464484
transform 1 0 36892 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1666464484
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_393
timestamp 1666464484
transform 1 0 37260 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_401
timestamp 1666464484
transform 1 0 37996 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_409
timestamp 1666464484
transform 1 0 38732 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_417
timestamp 1666464484
transform 1 0 39468 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_425
timestamp 1666464484
transform 1 0 40204 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_433
timestamp 1666464484
transform 1 0 40940 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_441
timestamp 1666464484
transform 1 0 41676 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_445
timestamp 1666464484
transform 1 0 42044 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1666464484
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_449
timestamp 1666464484
transform 1 0 42412 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_457
timestamp 1666464484
transform 1 0 43148 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_465
timestamp 1666464484
transform 1 0 43884 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_473
timestamp 1666464484
transform 1 0 44620 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_481
timestamp 1666464484
transform 1 0 45356 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_489
timestamp 1666464484
transform 1 0 46092 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_497
timestamp 1666464484
transform 1 0 46828 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_501
timestamp 1666464484
transform 1 0 47196 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1666464484
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_505
timestamp 1666464484
transform 1 0 47564 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_513
timestamp 1666464484
transform 1 0 48300 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_521
timestamp 1666464484
transform 1 0 49036 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_529
timestamp 1666464484
transform 1 0 49772 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_537
timestamp 1666464484
transform 1 0 50508 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_545
timestamp 1666464484
transform 1 0 51244 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_553
timestamp 1666464484
transform 1 0 51980 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_557
timestamp 1666464484
transform 1 0 52348 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1666464484
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_561
timestamp 1666464484
transform 1 0 52716 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_569
timestamp 1666464484
transform 1 0 53452 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_577
timestamp 1666464484
transform 1 0 54188 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_585
timestamp 1666464484
transform 1 0 54924 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_593
timestamp 1666464484
transform 1 0 55660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_79_601
timestamp 1666464484
transform 1 0 56396 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_79_609
timestamp 1666464484
transform 1 0 57132 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_613
timestamp 1666464484
transform 1 0 57500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1666464484
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_79_617
timestamp 1666464484
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_3
timestamp 1666464484
transform 1 0 1380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_11
timestamp 1666464484
transform 1 0 2116 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_19
timestamp 1666464484
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1666464484
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_29
timestamp 1666464484
transform 1 0 3772 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_37
timestamp 1666464484
transform 1 0 4508 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_45
timestamp 1666464484
transform 1 0 5244 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_53
timestamp 1666464484
transform 1 0 5980 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_61
timestamp 1666464484
transform 1 0 6716 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_69
timestamp 1666464484
transform 1 0 7452 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_77
timestamp 1666464484
transform 1 0 8188 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_81
timestamp 1666464484
transform 1 0 8556 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1666464484
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_85
timestamp 1666464484
transform 1 0 8924 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_93
timestamp 1666464484
transform 1 0 9660 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_101
timestamp 1666464484
transform 1 0 10396 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_109
timestamp 1666464484
transform 1 0 11132 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_117
timestamp 1666464484
transform 1 0 11868 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_125
timestamp 1666464484
transform 1 0 12604 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_133
timestamp 1666464484
transform 1 0 13340 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_137
timestamp 1666464484
transform 1 0 13708 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1666464484
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_141
timestamp 1666464484
transform 1 0 14076 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_149
timestamp 1666464484
transform 1 0 14812 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_157
timestamp 1666464484
transform 1 0 15548 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_165
timestamp 1666464484
transform 1 0 16284 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_173
timestamp 1666464484
transform 1 0 17020 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_181
timestamp 1666464484
transform 1 0 17756 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_189
timestamp 1666464484
transform 1 0 18492 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_193
timestamp 1666464484
transform 1 0 18860 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1666464484
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_197
timestamp 1666464484
transform 1 0 19228 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_205
timestamp 1666464484
transform 1 0 19964 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_213
timestamp 1666464484
transform 1 0 20700 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_221
timestamp 1666464484
transform 1 0 21436 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_229
timestamp 1666464484
transform 1 0 22172 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_237
timestamp 1666464484
transform 1 0 22908 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_245
timestamp 1666464484
transform 1 0 23644 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_249
timestamp 1666464484
transform 1 0 24012 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1666464484
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_253
timestamp 1666464484
transform 1 0 24380 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_261
timestamp 1666464484
transform 1 0 25116 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_269
timestamp 1666464484
transform 1 0 25852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_277
timestamp 1666464484
transform 1 0 26588 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_285
timestamp 1666464484
transform 1 0 27324 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_293
timestamp 1666464484
transform 1 0 28060 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_301
timestamp 1666464484
transform 1 0 28796 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_305
timestamp 1666464484
transform 1 0 29164 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1666464484
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_309
timestamp 1666464484
transform 1 0 29532 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_317
timestamp 1666464484
transform 1 0 30268 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_325
timestamp 1666464484
transform 1 0 31004 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_333
timestamp 1666464484
transform 1 0 31740 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_341
timestamp 1666464484
transform 1 0 32476 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_349
timestamp 1666464484
transform 1 0 33212 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_357
timestamp 1666464484
transform 1 0 33948 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_361
timestamp 1666464484
transform 1 0 34316 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1666464484
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_365
timestamp 1666464484
transform 1 0 34684 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_373
timestamp 1666464484
transform 1 0 35420 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_381
timestamp 1666464484
transform 1 0 36156 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_389
timestamp 1666464484
transform 1 0 36892 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_397
timestamp 1666464484
transform 1 0 37628 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_405
timestamp 1666464484
transform 1 0 38364 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_413
timestamp 1666464484
transform 1 0 39100 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_417
timestamp 1666464484
transform 1 0 39468 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1666464484
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_421
timestamp 1666464484
transform 1 0 39836 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_429
timestamp 1666464484
transform 1 0 40572 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_437
timestamp 1666464484
transform 1 0 41308 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_445
timestamp 1666464484
transform 1 0 42044 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_453
timestamp 1666464484
transform 1 0 42780 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_461
timestamp 1666464484
transform 1 0 43516 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_469
timestamp 1666464484
transform 1 0 44252 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_473
timestamp 1666464484
transform 1 0 44620 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1666464484
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_477
timestamp 1666464484
transform 1 0 44988 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_485
timestamp 1666464484
transform 1 0 45724 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_493
timestamp 1666464484
transform 1 0 46460 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_501
timestamp 1666464484
transform 1 0 47196 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_509
timestamp 1666464484
transform 1 0 47932 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_517
timestamp 1666464484
transform 1 0 48668 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_525
timestamp 1666464484
transform 1 0 49404 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_529
timestamp 1666464484
transform 1 0 49772 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1666464484
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_533
timestamp 1666464484
transform 1 0 50140 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_541
timestamp 1666464484
transform 1 0 50876 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_549
timestamp 1666464484
transform 1 0 51612 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_557
timestamp 1666464484
transform 1 0 52348 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_565
timestamp 1666464484
transform 1 0 53084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_573
timestamp 1666464484
transform 1 0 53820 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_581
timestamp 1666464484
transform 1 0 54556 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_585
timestamp 1666464484
transform 1 0 54924 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1666464484
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_80_589
timestamp 1666464484
transform 1 0 55292 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_597
timestamp 1666464484
transform 1 0 56028 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_605
timestamp 1666464484
transform 1 0 56764 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_80_613
timestamp 1666464484
transform 1 0 57500 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_80_621
timestamp 1666464484
transform 1 0 58236 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_81_3
timestamp 1666464484
transform 1 0 1380 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_11
timestamp 1666464484
transform 1 0 2116 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_19
timestamp 1666464484
transform 1 0 2852 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_27
timestamp 1666464484
transform 1 0 3588 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_35
timestamp 1666464484
transform 1 0 4324 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_43
timestamp 1666464484
transform 1 0 5060 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_51
timestamp 1666464484
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1666464484
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_57
timestamp 1666464484
transform 1 0 6348 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_65
timestamp 1666464484
transform 1 0 7084 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_73
timestamp 1666464484
transform 1 0 7820 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_81
timestamp 1666464484
transform 1 0 8556 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_89
timestamp 1666464484
transform 1 0 9292 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_97
timestamp 1666464484
transform 1 0 10028 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_105
timestamp 1666464484
transform 1 0 10764 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_109
timestamp 1666464484
transform 1 0 11132 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1666464484
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_113
timestamp 1666464484
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_121
timestamp 1666464484
transform 1 0 12236 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_129
timestamp 1666464484
transform 1 0 12972 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_137
timestamp 1666464484
transform 1 0 13708 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_145
timestamp 1666464484
transform 1 0 14444 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_153
timestamp 1666464484
transform 1 0 15180 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_161
timestamp 1666464484
transform 1 0 15916 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_165
timestamp 1666464484
transform 1 0 16284 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1666464484
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_169
timestamp 1666464484
transform 1 0 16652 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_177
timestamp 1666464484
transform 1 0 17388 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_185
timestamp 1666464484
transform 1 0 18124 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_193
timestamp 1666464484
transform 1 0 18860 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_201
timestamp 1666464484
transform 1 0 19596 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_209
timestamp 1666464484
transform 1 0 20332 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_217
timestamp 1666464484
transform 1 0 21068 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_221
timestamp 1666464484
transform 1 0 21436 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1666464484
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_225
timestamp 1666464484
transform 1 0 21804 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_233
timestamp 1666464484
transform 1 0 22540 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_241
timestamp 1666464484
transform 1 0 23276 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_249
timestamp 1666464484
transform 1 0 24012 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_257
timestamp 1666464484
transform 1 0 24748 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_265
timestamp 1666464484
transform 1 0 25484 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_273
timestamp 1666464484
transform 1 0 26220 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_277
timestamp 1666464484
transform 1 0 26588 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1666464484
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_281
timestamp 1666464484
transform 1 0 26956 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_289
timestamp 1666464484
transform 1 0 27692 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_297
timestamp 1666464484
transform 1 0 28428 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_305
timestamp 1666464484
transform 1 0 29164 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_313
timestamp 1666464484
transform 1 0 29900 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_321
timestamp 1666464484
transform 1 0 30636 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_329
timestamp 1666464484
transform 1 0 31372 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_333
timestamp 1666464484
transform 1 0 31740 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1666464484
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_337
timestamp 1666464484
transform 1 0 32108 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_345
timestamp 1666464484
transform 1 0 32844 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_353
timestamp 1666464484
transform 1 0 33580 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_361
timestamp 1666464484
transform 1 0 34316 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_369
timestamp 1666464484
transform 1 0 35052 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_377
timestamp 1666464484
transform 1 0 35788 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_385
timestamp 1666464484
transform 1 0 36524 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_389
timestamp 1666464484
transform 1 0 36892 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1666464484
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_393
timestamp 1666464484
transform 1 0 37260 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_401
timestamp 1666464484
transform 1 0 37996 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_409
timestamp 1666464484
transform 1 0 38732 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_417
timestamp 1666464484
transform 1 0 39468 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_425
timestamp 1666464484
transform 1 0 40204 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_433
timestamp 1666464484
transform 1 0 40940 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_441
timestamp 1666464484
transform 1 0 41676 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_445
timestamp 1666464484
transform 1 0 42044 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1666464484
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_449
timestamp 1666464484
transform 1 0 42412 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_457
timestamp 1666464484
transform 1 0 43148 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_465
timestamp 1666464484
transform 1 0 43884 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_473
timestamp 1666464484
transform 1 0 44620 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_481
timestamp 1666464484
transform 1 0 45356 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_489
timestamp 1666464484
transform 1 0 46092 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_497
timestamp 1666464484
transform 1 0 46828 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_501
timestamp 1666464484
transform 1 0 47196 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1666464484
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_505
timestamp 1666464484
transform 1 0 47564 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_513
timestamp 1666464484
transform 1 0 48300 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_521
timestamp 1666464484
transform 1 0 49036 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_529
timestamp 1666464484
transform 1 0 49772 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_537
timestamp 1666464484
transform 1 0 50508 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_545
timestamp 1666464484
transform 1 0 51244 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_553
timestamp 1666464484
transform 1 0 51980 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_557
timestamp 1666464484
transform 1 0 52348 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1666464484
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_561
timestamp 1666464484
transform 1 0 52716 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_569
timestamp 1666464484
transform 1 0 53452 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_577
timestamp 1666464484
transform 1 0 54188 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_585
timestamp 1666464484
transform 1 0 54924 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_593
timestamp 1666464484
transform 1 0 55660 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_81_601
timestamp 1666464484
transform 1 0 56396 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_81_609
timestamp 1666464484
transform 1 0 57132 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_613
timestamp 1666464484
transform 1 0 57500 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1666464484
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_81_617
timestamp 1666464484
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_3
timestamp 1666464484
transform 1 0 1380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_11
timestamp 1666464484
transform 1 0 2116 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_19
timestamp 1666464484
transform 1 0 2852 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1666464484
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_29
timestamp 1666464484
transform 1 0 3772 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_37
timestamp 1666464484
transform 1 0 4508 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_45
timestamp 1666464484
transform 1 0 5244 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_53
timestamp 1666464484
transform 1 0 5980 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_61
timestamp 1666464484
transform 1 0 6716 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_69
timestamp 1666464484
transform 1 0 7452 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_77
timestamp 1666464484
transform 1 0 8188 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_81
timestamp 1666464484
transform 1 0 8556 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1666464484
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_85
timestamp 1666464484
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_93
timestamp 1666464484
transform 1 0 9660 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_101
timestamp 1666464484
transform 1 0 10396 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_109
timestamp 1666464484
transform 1 0 11132 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_117
timestamp 1666464484
transform 1 0 11868 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_125
timestamp 1666464484
transform 1 0 12604 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_133
timestamp 1666464484
transform 1 0 13340 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_137
timestamp 1666464484
transform 1 0 13708 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1666464484
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_141
timestamp 1666464484
transform 1 0 14076 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_149
timestamp 1666464484
transform 1 0 14812 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_157
timestamp 1666464484
transform 1 0 15548 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_165
timestamp 1666464484
transform 1 0 16284 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_173
timestamp 1666464484
transform 1 0 17020 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_181
timestamp 1666464484
transform 1 0 17756 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_189
timestamp 1666464484
transform 1 0 18492 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_193
timestamp 1666464484
transform 1 0 18860 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1666464484
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_197
timestamp 1666464484
transform 1 0 19228 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_205
timestamp 1666464484
transform 1 0 19964 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_213
timestamp 1666464484
transform 1 0 20700 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_221
timestamp 1666464484
transform 1 0 21436 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_229
timestamp 1666464484
transform 1 0 22172 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_237
timestamp 1666464484
transform 1 0 22908 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_245
timestamp 1666464484
transform 1 0 23644 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_249
timestamp 1666464484
transform 1 0 24012 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1666464484
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_253
timestamp 1666464484
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_261
timestamp 1666464484
transform 1 0 25116 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_269
timestamp 1666464484
transform 1 0 25852 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_277
timestamp 1666464484
transform 1 0 26588 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_285
timestamp 1666464484
transform 1 0 27324 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_293
timestamp 1666464484
transform 1 0 28060 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_301
timestamp 1666464484
transform 1 0 28796 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_305
timestamp 1666464484
transform 1 0 29164 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1666464484
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_309
timestamp 1666464484
transform 1 0 29532 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_317
timestamp 1666464484
transform 1 0 30268 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_325
timestamp 1666464484
transform 1 0 31004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_333
timestamp 1666464484
transform 1 0 31740 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_341
timestamp 1666464484
transform 1 0 32476 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_349
timestamp 1666464484
transform 1 0 33212 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_357
timestamp 1666464484
transform 1 0 33948 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_361
timestamp 1666464484
transform 1 0 34316 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1666464484
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_365
timestamp 1666464484
transform 1 0 34684 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_373
timestamp 1666464484
transform 1 0 35420 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_381
timestamp 1666464484
transform 1 0 36156 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_389
timestamp 1666464484
transform 1 0 36892 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_397
timestamp 1666464484
transform 1 0 37628 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_405
timestamp 1666464484
transform 1 0 38364 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_413
timestamp 1666464484
transform 1 0 39100 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_417
timestamp 1666464484
transform 1 0 39468 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1666464484
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_421
timestamp 1666464484
transform 1 0 39836 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_429
timestamp 1666464484
transform 1 0 40572 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_437
timestamp 1666464484
transform 1 0 41308 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_445
timestamp 1666464484
transform 1 0 42044 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_453
timestamp 1666464484
transform 1 0 42780 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_461
timestamp 1666464484
transform 1 0 43516 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_469
timestamp 1666464484
transform 1 0 44252 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_473
timestamp 1666464484
transform 1 0 44620 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1666464484
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_477
timestamp 1666464484
transform 1 0 44988 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_485
timestamp 1666464484
transform 1 0 45724 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_493
timestamp 1666464484
transform 1 0 46460 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_501
timestamp 1666464484
transform 1 0 47196 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_509
timestamp 1666464484
transform 1 0 47932 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_517
timestamp 1666464484
transform 1 0 48668 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_525
timestamp 1666464484
transform 1 0 49404 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_529
timestamp 1666464484
transform 1 0 49772 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1666464484
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_533
timestamp 1666464484
transform 1 0 50140 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_541
timestamp 1666464484
transform 1 0 50876 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_549
timestamp 1666464484
transform 1 0 51612 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_557
timestamp 1666464484
transform 1 0 52348 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_565
timestamp 1666464484
transform 1 0 53084 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_573
timestamp 1666464484
transform 1 0 53820 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_581
timestamp 1666464484
transform 1 0 54556 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_585
timestamp 1666464484
transform 1 0 54924 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1666464484
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_82_589
timestamp 1666464484
transform 1 0 55292 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_597
timestamp 1666464484
transform 1 0 56028 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_605
timestamp 1666464484
transform 1 0 56764 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_82_613
timestamp 1666464484
transform 1 0 57500 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_82_621
timestamp 1666464484
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_83_3
timestamp 1666464484
transform 1 0 1380 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_11
timestamp 1666464484
transform 1 0 2116 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_19
timestamp 1666464484
transform 1 0 2852 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_27
timestamp 1666464484
transform 1 0 3588 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_35
timestamp 1666464484
transform 1 0 4324 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_43
timestamp 1666464484
transform 1 0 5060 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_51
timestamp 1666464484
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1666464484
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_57
timestamp 1666464484
transform 1 0 6348 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_65
timestamp 1666464484
transform 1 0 7084 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_73
timestamp 1666464484
transform 1 0 7820 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_81
timestamp 1666464484
transform 1 0 8556 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_89
timestamp 1666464484
transform 1 0 9292 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_97
timestamp 1666464484
transform 1 0 10028 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_105
timestamp 1666464484
transform 1 0 10764 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_109
timestamp 1666464484
transform 1 0 11132 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1666464484
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_113
timestamp 1666464484
transform 1 0 11500 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_121
timestamp 1666464484
transform 1 0 12236 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_129
timestamp 1666464484
transform 1 0 12972 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_137
timestamp 1666464484
transform 1 0 13708 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_145
timestamp 1666464484
transform 1 0 14444 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_153
timestamp 1666464484
transform 1 0 15180 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_161
timestamp 1666464484
transform 1 0 15916 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_165
timestamp 1666464484
transform 1 0 16284 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1666464484
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_169
timestamp 1666464484
transform 1 0 16652 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_177
timestamp 1666464484
transform 1 0 17388 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_185
timestamp 1666464484
transform 1 0 18124 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_193
timestamp 1666464484
transform 1 0 18860 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_201
timestamp 1666464484
transform 1 0 19596 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_209
timestamp 1666464484
transform 1 0 20332 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_217
timestamp 1666464484
transform 1 0 21068 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_221
timestamp 1666464484
transform 1 0 21436 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1666464484
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_225
timestamp 1666464484
transform 1 0 21804 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_233
timestamp 1666464484
transform 1 0 22540 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_241
timestamp 1666464484
transform 1 0 23276 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_249
timestamp 1666464484
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_257
timestamp 1666464484
transform 1 0 24748 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_265
timestamp 1666464484
transform 1 0 25484 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_273
timestamp 1666464484
transform 1 0 26220 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_277
timestamp 1666464484
transform 1 0 26588 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1666464484
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_281
timestamp 1666464484
transform 1 0 26956 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_289
timestamp 1666464484
transform 1 0 27692 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_297
timestamp 1666464484
transform 1 0 28428 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_305
timestamp 1666464484
transform 1 0 29164 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_313
timestamp 1666464484
transform 1 0 29900 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_321
timestamp 1666464484
transform 1 0 30636 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_329
timestamp 1666464484
transform 1 0 31372 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_333
timestamp 1666464484
transform 1 0 31740 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1666464484
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_337
timestamp 1666464484
transform 1 0 32108 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_345
timestamp 1666464484
transform 1 0 32844 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_353
timestamp 1666464484
transform 1 0 33580 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_361
timestamp 1666464484
transform 1 0 34316 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_369
timestamp 1666464484
transform 1 0 35052 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_377
timestamp 1666464484
transform 1 0 35788 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_385
timestamp 1666464484
transform 1 0 36524 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_389
timestamp 1666464484
transform 1 0 36892 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1666464484
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_393
timestamp 1666464484
transform 1 0 37260 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_401
timestamp 1666464484
transform 1 0 37996 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_409
timestamp 1666464484
transform 1 0 38732 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_417
timestamp 1666464484
transform 1 0 39468 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_425
timestamp 1666464484
transform 1 0 40204 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_433
timestamp 1666464484
transform 1 0 40940 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_441
timestamp 1666464484
transform 1 0 41676 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_445
timestamp 1666464484
transform 1 0 42044 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1666464484
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_449
timestamp 1666464484
transform 1 0 42412 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_457
timestamp 1666464484
transform 1 0 43148 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_465
timestamp 1666464484
transform 1 0 43884 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_473
timestamp 1666464484
transform 1 0 44620 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_481
timestamp 1666464484
transform 1 0 45356 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_489
timestamp 1666464484
transform 1 0 46092 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_497
timestamp 1666464484
transform 1 0 46828 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_501
timestamp 1666464484
transform 1 0 47196 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1666464484
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_505
timestamp 1666464484
transform 1 0 47564 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_513
timestamp 1666464484
transform 1 0 48300 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_521
timestamp 1666464484
transform 1 0 49036 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_529
timestamp 1666464484
transform 1 0 49772 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_537
timestamp 1666464484
transform 1 0 50508 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_545
timestamp 1666464484
transform 1 0 51244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_553
timestamp 1666464484
transform 1 0 51980 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_557
timestamp 1666464484
transform 1 0 52348 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1666464484
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_561
timestamp 1666464484
transform 1 0 52716 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_569
timestamp 1666464484
transform 1 0 53452 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_577
timestamp 1666464484
transform 1 0 54188 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_585
timestamp 1666464484
transform 1 0 54924 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_593
timestamp 1666464484
transform 1 0 55660 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_83_601
timestamp 1666464484
transform 1 0 56396 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_83_609
timestamp 1666464484
transform 1 0 57132 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_613
timestamp 1666464484
transform 1 0 57500 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1666464484
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_83_617
timestamp 1666464484
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_3
timestamp 1666464484
transform 1 0 1380 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_11
timestamp 1666464484
transform 1 0 2116 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_19
timestamp 1666464484
transform 1 0 2852 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1666464484
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_29
timestamp 1666464484
transform 1 0 3772 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_37
timestamp 1666464484
transform 1 0 4508 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_45
timestamp 1666464484
transform 1 0 5244 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_53
timestamp 1666464484
transform 1 0 5980 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_61
timestamp 1666464484
transform 1 0 6716 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_69
timestamp 1666464484
transform 1 0 7452 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_77
timestamp 1666464484
transform 1 0 8188 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_81
timestamp 1666464484
transform 1 0 8556 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1666464484
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_85
timestamp 1666464484
transform 1 0 8924 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_93
timestamp 1666464484
transform 1 0 9660 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_101
timestamp 1666464484
transform 1 0 10396 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_109
timestamp 1666464484
transform 1 0 11132 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_117
timestamp 1666464484
transform 1 0 11868 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_125
timestamp 1666464484
transform 1 0 12604 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_133
timestamp 1666464484
transform 1 0 13340 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_137
timestamp 1666464484
transform 1 0 13708 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1666464484
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_141
timestamp 1666464484
transform 1 0 14076 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_149
timestamp 1666464484
transform 1 0 14812 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_157
timestamp 1666464484
transform 1 0 15548 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_165
timestamp 1666464484
transform 1 0 16284 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_173
timestamp 1666464484
transform 1 0 17020 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_181
timestamp 1666464484
transform 1 0 17756 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_189
timestamp 1666464484
transform 1 0 18492 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_193
timestamp 1666464484
transform 1 0 18860 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1666464484
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_197
timestamp 1666464484
transform 1 0 19228 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_205
timestamp 1666464484
transform 1 0 19964 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_213
timestamp 1666464484
transform 1 0 20700 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_221
timestamp 1666464484
transform 1 0 21436 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_229
timestamp 1666464484
transform 1 0 22172 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_237
timestamp 1666464484
transform 1 0 22908 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_245
timestamp 1666464484
transform 1 0 23644 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_249
timestamp 1666464484
transform 1 0 24012 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1666464484
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_253
timestamp 1666464484
transform 1 0 24380 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_261
timestamp 1666464484
transform 1 0 25116 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_269
timestamp 1666464484
transform 1 0 25852 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_277
timestamp 1666464484
transform 1 0 26588 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_285
timestamp 1666464484
transform 1 0 27324 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_293
timestamp 1666464484
transform 1 0 28060 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_301
timestamp 1666464484
transform 1 0 28796 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_305
timestamp 1666464484
transform 1 0 29164 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1666464484
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_309
timestamp 1666464484
transform 1 0 29532 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_317
timestamp 1666464484
transform 1 0 30268 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_325
timestamp 1666464484
transform 1 0 31004 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_333
timestamp 1666464484
transform 1 0 31740 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_341
timestamp 1666464484
transform 1 0 32476 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_349
timestamp 1666464484
transform 1 0 33212 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_357
timestamp 1666464484
transform 1 0 33948 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_361
timestamp 1666464484
transform 1 0 34316 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1666464484
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_365
timestamp 1666464484
transform 1 0 34684 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_373
timestamp 1666464484
transform 1 0 35420 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_381
timestamp 1666464484
transform 1 0 36156 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_389
timestamp 1666464484
transform 1 0 36892 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_397
timestamp 1666464484
transform 1 0 37628 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_405
timestamp 1666464484
transform 1 0 38364 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_413
timestamp 1666464484
transform 1 0 39100 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_417
timestamp 1666464484
transform 1 0 39468 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1666464484
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_421
timestamp 1666464484
transform 1 0 39836 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_429
timestamp 1666464484
transform 1 0 40572 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_437
timestamp 1666464484
transform 1 0 41308 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_445
timestamp 1666464484
transform 1 0 42044 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_453
timestamp 1666464484
transform 1 0 42780 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_461
timestamp 1666464484
transform 1 0 43516 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_469
timestamp 1666464484
transform 1 0 44252 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_473
timestamp 1666464484
transform 1 0 44620 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1666464484
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_477
timestamp 1666464484
transform 1 0 44988 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_485
timestamp 1666464484
transform 1 0 45724 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_493
timestamp 1666464484
transform 1 0 46460 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_501
timestamp 1666464484
transform 1 0 47196 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_509
timestamp 1666464484
transform 1 0 47932 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_517
timestamp 1666464484
transform 1 0 48668 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_525
timestamp 1666464484
transform 1 0 49404 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_529
timestamp 1666464484
transform 1 0 49772 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1666464484
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_533
timestamp 1666464484
transform 1 0 50140 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_541
timestamp 1666464484
transform 1 0 50876 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_549
timestamp 1666464484
transform 1 0 51612 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_557
timestamp 1666464484
transform 1 0 52348 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_565
timestamp 1666464484
transform 1 0 53084 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_573
timestamp 1666464484
transform 1 0 53820 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_581
timestamp 1666464484
transform 1 0 54556 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_585
timestamp 1666464484
transform 1 0 54924 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1666464484
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_84_589
timestamp 1666464484
transform 1 0 55292 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_597
timestamp 1666464484
transform 1 0 56028 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_605
timestamp 1666464484
transform 1 0 56764 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_84_613
timestamp 1666464484
transform 1 0 57500 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_84_621
timestamp 1666464484
transform 1 0 58236 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_85_3
timestamp 1666464484
transform 1 0 1380 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_11
timestamp 1666464484
transform 1 0 2116 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_19
timestamp 1666464484
transform 1 0 2852 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_27
timestamp 1666464484
transform 1 0 3588 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_35
timestamp 1666464484
transform 1 0 4324 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_43
timestamp 1666464484
transform 1 0 5060 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_51
timestamp 1666464484
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1666464484
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_57
timestamp 1666464484
transform 1 0 6348 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_65
timestamp 1666464484
transform 1 0 7084 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_73
timestamp 1666464484
transform 1 0 7820 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_81
timestamp 1666464484
transform 1 0 8556 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_89
timestamp 1666464484
transform 1 0 9292 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_97
timestamp 1666464484
transform 1 0 10028 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_105
timestamp 1666464484
transform 1 0 10764 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_109
timestamp 1666464484
transform 1 0 11132 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1666464484
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_113
timestamp 1666464484
transform 1 0 11500 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_121
timestamp 1666464484
transform 1 0 12236 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_129
timestamp 1666464484
transform 1 0 12972 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_137
timestamp 1666464484
transform 1 0 13708 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_145
timestamp 1666464484
transform 1 0 14444 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_153
timestamp 1666464484
transform 1 0 15180 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_161
timestamp 1666464484
transform 1 0 15916 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_165
timestamp 1666464484
transform 1 0 16284 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1666464484
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_169
timestamp 1666464484
transform 1 0 16652 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_177
timestamp 1666464484
transform 1 0 17388 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_185
timestamp 1666464484
transform 1 0 18124 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_193
timestamp 1666464484
transform 1 0 18860 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_201
timestamp 1666464484
transform 1 0 19596 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_209
timestamp 1666464484
transform 1 0 20332 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_217
timestamp 1666464484
transform 1 0 21068 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_221
timestamp 1666464484
transform 1 0 21436 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1666464484
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_225
timestamp 1666464484
transform 1 0 21804 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_233
timestamp 1666464484
transform 1 0 22540 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_241
timestamp 1666464484
transform 1 0 23276 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_249
timestamp 1666464484
transform 1 0 24012 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_257
timestamp 1666464484
transform 1 0 24748 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_265
timestamp 1666464484
transform 1 0 25484 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_273
timestamp 1666464484
transform 1 0 26220 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_277
timestamp 1666464484
transform 1 0 26588 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1666464484
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_281
timestamp 1666464484
transform 1 0 26956 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_289
timestamp 1666464484
transform 1 0 27692 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_297
timestamp 1666464484
transform 1 0 28428 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_305
timestamp 1666464484
transform 1 0 29164 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_313
timestamp 1666464484
transform 1 0 29900 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_321
timestamp 1666464484
transform 1 0 30636 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_329
timestamp 1666464484
transform 1 0 31372 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_333
timestamp 1666464484
transform 1 0 31740 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1666464484
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_337
timestamp 1666464484
transform 1 0 32108 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_345
timestamp 1666464484
transform 1 0 32844 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_353
timestamp 1666464484
transform 1 0 33580 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_361
timestamp 1666464484
transform 1 0 34316 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_369
timestamp 1666464484
transform 1 0 35052 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_377
timestamp 1666464484
transform 1 0 35788 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_385
timestamp 1666464484
transform 1 0 36524 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_389
timestamp 1666464484
transform 1 0 36892 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1666464484
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_393
timestamp 1666464484
transform 1 0 37260 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_401
timestamp 1666464484
transform 1 0 37996 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_409
timestamp 1666464484
transform 1 0 38732 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_417
timestamp 1666464484
transform 1 0 39468 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_425
timestamp 1666464484
transform 1 0 40204 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_433
timestamp 1666464484
transform 1 0 40940 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_441
timestamp 1666464484
transform 1 0 41676 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_445
timestamp 1666464484
transform 1 0 42044 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1666464484
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_449
timestamp 1666464484
transform 1 0 42412 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_457
timestamp 1666464484
transform 1 0 43148 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_465
timestamp 1666464484
transform 1 0 43884 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_473
timestamp 1666464484
transform 1 0 44620 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_481
timestamp 1666464484
transform 1 0 45356 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_489
timestamp 1666464484
transform 1 0 46092 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_497
timestamp 1666464484
transform 1 0 46828 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_501
timestamp 1666464484
transform 1 0 47196 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1666464484
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_505
timestamp 1666464484
transform 1 0 47564 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_513
timestamp 1666464484
transform 1 0 48300 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_521
timestamp 1666464484
transform 1 0 49036 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_529
timestamp 1666464484
transform 1 0 49772 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_537
timestamp 1666464484
transform 1 0 50508 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_545
timestamp 1666464484
transform 1 0 51244 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_553
timestamp 1666464484
transform 1 0 51980 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_557
timestamp 1666464484
transform 1 0 52348 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1666464484
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_561
timestamp 1666464484
transform 1 0 52716 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_569
timestamp 1666464484
transform 1 0 53452 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_577
timestamp 1666464484
transform 1 0 54188 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_585
timestamp 1666464484
transform 1 0 54924 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_593
timestamp 1666464484
transform 1 0 55660 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_85_601
timestamp 1666464484
transform 1 0 56396 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_85_609
timestamp 1666464484
transform 1 0 57132 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_613
timestamp 1666464484
transform 1 0 57500 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1666464484
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_85_617
timestamp 1666464484
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_3
timestamp 1666464484
transform 1 0 1380 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_11
timestamp 1666464484
transform 1 0 2116 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_19
timestamp 1666464484
transform 1 0 2852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1666464484
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_29
timestamp 1666464484
transform 1 0 3772 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_37
timestamp 1666464484
transform 1 0 4508 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_45
timestamp 1666464484
transform 1 0 5244 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_53
timestamp 1666464484
transform 1 0 5980 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_61
timestamp 1666464484
transform 1 0 6716 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_69
timestamp 1666464484
transform 1 0 7452 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_77
timestamp 1666464484
transform 1 0 8188 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_81
timestamp 1666464484
transform 1 0 8556 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1666464484
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_85
timestamp 1666464484
transform 1 0 8924 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_93
timestamp 1666464484
transform 1 0 9660 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_101
timestamp 1666464484
transform 1 0 10396 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_109
timestamp 1666464484
transform 1 0 11132 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_117
timestamp 1666464484
transform 1 0 11868 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_125
timestamp 1666464484
transform 1 0 12604 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_133
timestamp 1666464484
transform 1 0 13340 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_137
timestamp 1666464484
transform 1 0 13708 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1666464484
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_141
timestamp 1666464484
transform 1 0 14076 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_149
timestamp 1666464484
transform 1 0 14812 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_157
timestamp 1666464484
transform 1 0 15548 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_165
timestamp 1666464484
transform 1 0 16284 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_173
timestamp 1666464484
transform 1 0 17020 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_181
timestamp 1666464484
transform 1 0 17756 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_189
timestamp 1666464484
transform 1 0 18492 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_193
timestamp 1666464484
transform 1 0 18860 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1666464484
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_197
timestamp 1666464484
transform 1 0 19228 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_205
timestamp 1666464484
transform 1 0 19964 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_213
timestamp 1666464484
transform 1 0 20700 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_221
timestamp 1666464484
transform 1 0 21436 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_229
timestamp 1666464484
transform 1 0 22172 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_237
timestamp 1666464484
transform 1 0 22908 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_245
timestamp 1666464484
transform 1 0 23644 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_249
timestamp 1666464484
transform 1 0 24012 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1666464484
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_253
timestamp 1666464484
transform 1 0 24380 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_261
timestamp 1666464484
transform 1 0 25116 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_269
timestamp 1666464484
transform 1 0 25852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_277
timestamp 1666464484
transform 1 0 26588 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_285
timestamp 1666464484
transform 1 0 27324 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_293
timestamp 1666464484
transform 1 0 28060 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_301
timestamp 1666464484
transform 1 0 28796 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_305
timestamp 1666464484
transform 1 0 29164 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1666464484
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_309
timestamp 1666464484
transform 1 0 29532 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_317
timestamp 1666464484
transform 1 0 30268 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_325
timestamp 1666464484
transform 1 0 31004 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_333
timestamp 1666464484
transform 1 0 31740 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_341
timestamp 1666464484
transform 1 0 32476 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_349
timestamp 1666464484
transform 1 0 33212 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_357
timestamp 1666464484
transform 1 0 33948 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_361
timestamp 1666464484
transform 1 0 34316 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1666464484
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_365
timestamp 1666464484
transform 1 0 34684 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_373
timestamp 1666464484
transform 1 0 35420 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_381
timestamp 1666464484
transform 1 0 36156 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_389
timestamp 1666464484
transform 1 0 36892 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_397
timestamp 1666464484
transform 1 0 37628 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_405
timestamp 1666464484
transform 1 0 38364 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_413
timestamp 1666464484
transform 1 0 39100 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_417
timestamp 1666464484
transform 1 0 39468 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1666464484
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_421
timestamp 1666464484
transform 1 0 39836 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_429
timestamp 1666464484
transform 1 0 40572 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_437
timestamp 1666464484
transform 1 0 41308 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_445
timestamp 1666464484
transform 1 0 42044 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_453
timestamp 1666464484
transform 1 0 42780 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_461
timestamp 1666464484
transform 1 0 43516 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_469
timestamp 1666464484
transform 1 0 44252 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_473
timestamp 1666464484
transform 1 0 44620 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1666464484
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_477
timestamp 1666464484
transform 1 0 44988 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_485
timestamp 1666464484
transform 1 0 45724 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_493
timestamp 1666464484
transform 1 0 46460 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_501
timestamp 1666464484
transform 1 0 47196 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_509
timestamp 1666464484
transform 1 0 47932 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_517
timestamp 1666464484
transform 1 0 48668 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_525
timestamp 1666464484
transform 1 0 49404 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_529
timestamp 1666464484
transform 1 0 49772 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1666464484
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_533
timestamp 1666464484
transform 1 0 50140 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_541
timestamp 1666464484
transform 1 0 50876 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_549
timestamp 1666464484
transform 1 0 51612 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_557
timestamp 1666464484
transform 1 0 52348 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_565
timestamp 1666464484
transform 1 0 53084 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_573
timestamp 1666464484
transform 1 0 53820 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_581
timestamp 1666464484
transform 1 0 54556 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_585
timestamp 1666464484
transform 1 0 54924 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1666464484
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_86_589
timestamp 1666464484
transform 1 0 55292 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_597
timestamp 1666464484
transform 1 0 56028 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_605
timestamp 1666464484
transform 1 0 56764 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_86_613
timestamp 1666464484
transform 1 0 57500 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_86_621
timestamp 1666464484
transform 1 0 58236 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_87_3
timestamp 1666464484
transform 1 0 1380 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_11
timestamp 1666464484
transform 1 0 2116 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_19
timestamp 1666464484
transform 1 0 2852 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_27
timestamp 1666464484
transform 1 0 3588 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_35
timestamp 1666464484
transform 1 0 4324 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_43
timestamp 1666464484
transform 1 0 5060 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_51
timestamp 1666464484
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1666464484
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_57
timestamp 1666464484
transform 1 0 6348 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_65
timestamp 1666464484
transform 1 0 7084 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_73
timestamp 1666464484
transform 1 0 7820 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_81
timestamp 1666464484
transform 1 0 8556 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_89
timestamp 1666464484
transform 1 0 9292 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_97
timestamp 1666464484
transform 1 0 10028 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_105
timestamp 1666464484
transform 1 0 10764 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_109
timestamp 1666464484
transform 1 0 11132 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1666464484
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_113
timestamp 1666464484
transform 1 0 11500 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_121
timestamp 1666464484
transform 1 0 12236 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_129
timestamp 1666464484
transform 1 0 12972 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_137
timestamp 1666464484
transform 1 0 13708 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_145
timestamp 1666464484
transform 1 0 14444 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_153
timestamp 1666464484
transform 1 0 15180 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_161
timestamp 1666464484
transform 1 0 15916 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_165
timestamp 1666464484
transform 1 0 16284 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1666464484
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_169
timestamp 1666464484
transform 1 0 16652 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_177
timestamp 1666464484
transform 1 0 17388 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_185
timestamp 1666464484
transform 1 0 18124 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_193
timestamp 1666464484
transform 1 0 18860 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_201
timestamp 1666464484
transform 1 0 19596 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_209
timestamp 1666464484
transform 1 0 20332 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_217
timestamp 1666464484
transform 1 0 21068 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_221
timestamp 1666464484
transform 1 0 21436 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1666464484
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_225
timestamp 1666464484
transform 1 0 21804 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_233
timestamp 1666464484
transform 1 0 22540 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_241
timestamp 1666464484
transform 1 0 23276 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_249
timestamp 1666464484
transform 1 0 24012 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_257
timestamp 1666464484
transform 1 0 24748 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_265
timestamp 1666464484
transform 1 0 25484 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_273
timestamp 1666464484
transform 1 0 26220 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_277
timestamp 1666464484
transform 1 0 26588 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1666464484
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_281
timestamp 1666464484
transform 1 0 26956 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_289
timestamp 1666464484
transform 1 0 27692 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_297
timestamp 1666464484
transform 1 0 28428 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_305
timestamp 1666464484
transform 1 0 29164 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_313
timestamp 1666464484
transform 1 0 29900 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_321
timestamp 1666464484
transform 1 0 30636 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_329
timestamp 1666464484
transform 1 0 31372 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_333
timestamp 1666464484
transform 1 0 31740 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1666464484
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_337
timestamp 1666464484
transform 1 0 32108 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_345
timestamp 1666464484
transform 1 0 32844 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_353
timestamp 1666464484
transform 1 0 33580 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_361
timestamp 1666464484
transform 1 0 34316 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_369
timestamp 1666464484
transform 1 0 35052 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_377
timestamp 1666464484
transform 1 0 35788 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_385
timestamp 1666464484
transform 1 0 36524 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_389
timestamp 1666464484
transform 1 0 36892 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1666464484
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_393
timestamp 1666464484
transform 1 0 37260 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_401
timestamp 1666464484
transform 1 0 37996 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_409
timestamp 1666464484
transform 1 0 38732 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_417
timestamp 1666464484
transform 1 0 39468 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_425
timestamp 1666464484
transform 1 0 40204 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_433
timestamp 1666464484
transform 1 0 40940 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_441
timestamp 1666464484
transform 1 0 41676 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_445
timestamp 1666464484
transform 1 0 42044 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1666464484
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_449
timestamp 1666464484
transform 1 0 42412 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_457
timestamp 1666464484
transform 1 0 43148 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_465
timestamp 1666464484
transform 1 0 43884 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_473
timestamp 1666464484
transform 1 0 44620 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_481
timestamp 1666464484
transform 1 0 45356 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_489
timestamp 1666464484
transform 1 0 46092 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_497
timestamp 1666464484
transform 1 0 46828 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_501
timestamp 1666464484
transform 1 0 47196 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1666464484
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_505
timestamp 1666464484
transform 1 0 47564 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_513
timestamp 1666464484
transform 1 0 48300 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_521
timestamp 1666464484
transform 1 0 49036 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_529
timestamp 1666464484
transform 1 0 49772 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_537
timestamp 1666464484
transform 1 0 50508 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_545
timestamp 1666464484
transform 1 0 51244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_553
timestamp 1666464484
transform 1 0 51980 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_557
timestamp 1666464484
transform 1 0 52348 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1666464484
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_561
timestamp 1666464484
transform 1 0 52716 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_569
timestamp 1666464484
transform 1 0 53452 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_577
timestamp 1666464484
transform 1 0 54188 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_585
timestamp 1666464484
transform 1 0 54924 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_593
timestamp 1666464484
transform 1 0 55660 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_87_601
timestamp 1666464484
transform 1 0 56396 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_87_609
timestamp 1666464484
transform 1 0 57132 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_613
timestamp 1666464484
transform 1 0 57500 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1666464484
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_87_617
timestamp 1666464484
transform 1 0 57868 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_3
timestamp 1666464484
transform 1 0 1380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_11
timestamp 1666464484
transform 1 0 2116 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_19
timestamp 1666464484
transform 1 0 2852 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1666464484
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_29
timestamp 1666464484
transform 1 0 3772 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_37
timestamp 1666464484
transform 1 0 4508 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_45
timestamp 1666464484
transform 1 0 5244 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_53
timestamp 1666464484
transform 1 0 5980 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_61
timestamp 1666464484
transform 1 0 6716 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_69
timestamp 1666464484
transform 1 0 7452 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_77
timestamp 1666464484
transform 1 0 8188 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_81
timestamp 1666464484
transform 1 0 8556 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1666464484
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_85
timestamp 1666464484
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_93
timestamp 1666464484
transform 1 0 9660 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_101
timestamp 1666464484
transform 1 0 10396 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_109
timestamp 1666464484
transform 1 0 11132 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_117
timestamp 1666464484
transform 1 0 11868 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_125
timestamp 1666464484
transform 1 0 12604 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_133
timestamp 1666464484
transform 1 0 13340 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_137
timestamp 1666464484
transform 1 0 13708 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1666464484
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_141
timestamp 1666464484
transform 1 0 14076 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_149
timestamp 1666464484
transform 1 0 14812 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_157
timestamp 1666464484
transform 1 0 15548 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_165
timestamp 1666464484
transform 1 0 16284 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_173
timestamp 1666464484
transform 1 0 17020 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_181
timestamp 1666464484
transform 1 0 17756 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_189
timestamp 1666464484
transform 1 0 18492 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_193
timestamp 1666464484
transform 1 0 18860 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1666464484
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_197
timestamp 1666464484
transform 1 0 19228 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_205
timestamp 1666464484
transform 1 0 19964 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_213
timestamp 1666464484
transform 1 0 20700 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_221
timestamp 1666464484
transform 1 0 21436 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_229
timestamp 1666464484
transform 1 0 22172 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_237
timestamp 1666464484
transform 1 0 22908 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_245
timestamp 1666464484
transform 1 0 23644 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_249
timestamp 1666464484
transform 1 0 24012 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1666464484
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_253
timestamp 1666464484
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_261
timestamp 1666464484
transform 1 0 25116 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_269
timestamp 1666464484
transform 1 0 25852 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_277
timestamp 1666464484
transform 1 0 26588 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_285
timestamp 1666464484
transform 1 0 27324 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_293
timestamp 1666464484
transform 1 0 28060 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_301
timestamp 1666464484
transform 1 0 28796 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_305
timestamp 1666464484
transform 1 0 29164 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1666464484
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_309
timestamp 1666464484
transform 1 0 29532 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_317
timestamp 1666464484
transform 1 0 30268 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_325
timestamp 1666464484
transform 1 0 31004 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_333
timestamp 1666464484
transform 1 0 31740 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_341
timestamp 1666464484
transform 1 0 32476 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_349
timestamp 1666464484
transform 1 0 33212 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_357
timestamp 1666464484
transform 1 0 33948 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_361
timestamp 1666464484
transform 1 0 34316 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1666464484
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_365
timestamp 1666464484
transform 1 0 34684 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_373
timestamp 1666464484
transform 1 0 35420 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_381
timestamp 1666464484
transform 1 0 36156 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_389
timestamp 1666464484
transform 1 0 36892 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_397
timestamp 1666464484
transform 1 0 37628 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_405
timestamp 1666464484
transform 1 0 38364 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_413
timestamp 1666464484
transform 1 0 39100 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_417
timestamp 1666464484
transform 1 0 39468 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1666464484
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_421
timestamp 1666464484
transform 1 0 39836 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_429
timestamp 1666464484
transform 1 0 40572 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_437
timestamp 1666464484
transform 1 0 41308 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_445
timestamp 1666464484
transform 1 0 42044 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_453
timestamp 1666464484
transform 1 0 42780 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_461
timestamp 1666464484
transform 1 0 43516 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_469
timestamp 1666464484
transform 1 0 44252 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_473
timestamp 1666464484
transform 1 0 44620 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1666464484
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_477
timestamp 1666464484
transform 1 0 44988 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_485
timestamp 1666464484
transform 1 0 45724 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_493
timestamp 1666464484
transform 1 0 46460 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_501
timestamp 1666464484
transform 1 0 47196 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_509
timestamp 1666464484
transform 1 0 47932 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_517
timestamp 1666464484
transform 1 0 48668 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_525
timestamp 1666464484
transform 1 0 49404 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_529
timestamp 1666464484
transform 1 0 49772 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1666464484
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_533
timestamp 1666464484
transform 1 0 50140 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_541
timestamp 1666464484
transform 1 0 50876 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_549
timestamp 1666464484
transform 1 0 51612 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_557
timestamp 1666464484
transform 1 0 52348 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_565
timestamp 1666464484
transform 1 0 53084 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_573
timestamp 1666464484
transform 1 0 53820 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_581
timestamp 1666464484
transform 1 0 54556 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_88_585
timestamp 1666464484
transform 1 0 54924 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1666464484
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_88_589
timestamp 1666464484
transform 1 0 55292 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_597
timestamp 1666464484
transform 1 0 56028 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_605
timestamp 1666464484
transform 1 0 56764 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_88_613
timestamp 1666464484
transform 1 0 57500 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_88_621
timestamp 1666464484
transform 1 0 58236 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_89_3
timestamp 1666464484
transform 1 0 1380 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_11
timestamp 1666464484
transform 1 0 2116 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_19
timestamp 1666464484
transform 1 0 2852 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_27
timestamp 1666464484
transform 1 0 3588 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_35
timestamp 1666464484
transform 1 0 4324 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_43
timestamp 1666464484
transform 1 0 5060 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_51
timestamp 1666464484
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1666464484
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_57
timestamp 1666464484
transform 1 0 6348 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_65
timestamp 1666464484
transform 1 0 7084 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_73
timestamp 1666464484
transform 1 0 7820 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_81
timestamp 1666464484
transform 1 0 8556 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_89
timestamp 1666464484
transform 1 0 9292 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_97
timestamp 1666464484
transform 1 0 10028 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_105
timestamp 1666464484
transform 1 0 10764 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_109
timestamp 1666464484
transform 1 0 11132 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1666464484
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_113
timestamp 1666464484
transform 1 0 11500 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_121
timestamp 1666464484
transform 1 0 12236 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_129
timestamp 1666464484
transform 1 0 12972 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_137
timestamp 1666464484
transform 1 0 13708 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_145
timestamp 1666464484
transform 1 0 14444 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_153
timestamp 1666464484
transform 1 0 15180 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_161
timestamp 1666464484
transform 1 0 15916 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_165
timestamp 1666464484
transform 1 0 16284 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1666464484
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_169
timestamp 1666464484
transform 1 0 16652 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_177
timestamp 1666464484
transform 1 0 17388 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_185
timestamp 1666464484
transform 1 0 18124 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_193
timestamp 1666464484
transform 1 0 18860 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_201
timestamp 1666464484
transform 1 0 19596 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_209
timestamp 1666464484
transform 1 0 20332 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_217
timestamp 1666464484
transform 1 0 21068 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_221
timestamp 1666464484
transform 1 0 21436 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1666464484
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_225
timestamp 1666464484
transform 1 0 21804 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_233
timestamp 1666464484
transform 1 0 22540 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_241
timestamp 1666464484
transform 1 0 23276 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_249
timestamp 1666464484
transform 1 0 24012 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_257
timestamp 1666464484
transform 1 0 24748 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_265
timestamp 1666464484
transform 1 0 25484 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_273
timestamp 1666464484
transform 1 0 26220 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_277
timestamp 1666464484
transform 1 0 26588 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1666464484
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_281
timestamp 1666464484
transform 1 0 26956 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_289
timestamp 1666464484
transform 1 0 27692 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_297
timestamp 1666464484
transform 1 0 28428 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_305
timestamp 1666464484
transform 1 0 29164 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_313
timestamp 1666464484
transform 1 0 29900 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_321
timestamp 1666464484
transform 1 0 30636 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_329
timestamp 1666464484
transform 1 0 31372 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_333
timestamp 1666464484
transform 1 0 31740 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1666464484
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_337
timestamp 1666464484
transform 1 0 32108 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_345
timestamp 1666464484
transform 1 0 32844 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_353
timestamp 1666464484
transform 1 0 33580 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_361
timestamp 1666464484
transform 1 0 34316 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_369
timestamp 1666464484
transform 1 0 35052 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_377
timestamp 1666464484
transform 1 0 35788 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_385
timestamp 1666464484
transform 1 0 36524 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_389
timestamp 1666464484
transform 1 0 36892 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1666464484
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_393
timestamp 1666464484
transform 1 0 37260 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_401
timestamp 1666464484
transform 1 0 37996 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_409
timestamp 1666464484
transform 1 0 38732 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_417
timestamp 1666464484
transform 1 0 39468 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_425
timestamp 1666464484
transform 1 0 40204 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_433
timestamp 1666464484
transform 1 0 40940 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_441
timestamp 1666464484
transform 1 0 41676 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_445
timestamp 1666464484
transform 1 0 42044 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1666464484
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_449
timestamp 1666464484
transform 1 0 42412 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_457
timestamp 1666464484
transform 1 0 43148 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_465
timestamp 1666464484
transform 1 0 43884 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_473
timestamp 1666464484
transform 1 0 44620 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_481
timestamp 1666464484
transform 1 0 45356 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_489
timestamp 1666464484
transform 1 0 46092 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_497
timestamp 1666464484
transform 1 0 46828 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_501
timestamp 1666464484
transform 1 0 47196 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1666464484
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_505
timestamp 1666464484
transform 1 0 47564 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_513
timestamp 1666464484
transform 1 0 48300 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_521
timestamp 1666464484
transform 1 0 49036 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_529
timestamp 1666464484
transform 1 0 49772 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_537
timestamp 1666464484
transform 1 0 50508 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_545
timestamp 1666464484
transform 1 0 51244 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_553
timestamp 1666464484
transform 1 0 51980 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_557
timestamp 1666464484
transform 1 0 52348 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1666464484
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_561
timestamp 1666464484
transform 1 0 52716 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_569
timestamp 1666464484
transform 1 0 53452 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_577
timestamp 1666464484
transform 1 0 54188 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_585
timestamp 1666464484
transform 1 0 54924 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_593
timestamp 1666464484
transform 1 0 55660 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_89_601
timestamp 1666464484
transform 1 0 56396 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_89_609
timestamp 1666464484
transform 1 0 57132 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_613
timestamp 1666464484
transform 1 0 57500 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1666464484
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_89_617
timestamp 1666464484
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_3
timestamp 1666464484
transform 1 0 1380 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_11
timestamp 1666464484
transform 1 0 2116 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_19
timestamp 1666464484
transform 1 0 2852 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1666464484
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_29
timestamp 1666464484
transform 1 0 3772 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_37
timestamp 1666464484
transform 1 0 4508 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_45
timestamp 1666464484
transform 1 0 5244 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_53
timestamp 1666464484
transform 1 0 5980 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_61
timestamp 1666464484
transform 1 0 6716 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_69
timestamp 1666464484
transform 1 0 7452 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_77
timestamp 1666464484
transform 1 0 8188 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_81
timestamp 1666464484
transform 1 0 8556 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1666464484
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_85
timestamp 1666464484
transform 1 0 8924 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_93
timestamp 1666464484
transform 1 0 9660 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_101
timestamp 1666464484
transform 1 0 10396 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_109
timestamp 1666464484
transform 1 0 11132 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_117
timestamp 1666464484
transform 1 0 11868 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_125
timestamp 1666464484
transform 1 0 12604 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_133
timestamp 1666464484
transform 1 0 13340 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_137
timestamp 1666464484
transform 1 0 13708 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1666464484
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_141
timestamp 1666464484
transform 1 0 14076 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_149
timestamp 1666464484
transform 1 0 14812 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_157
timestamp 1666464484
transform 1 0 15548 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_165
timestamp 1666464484
transform 1 0 16284 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_173
timestamp 1666464484
transform 1 0 17020 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_181
timestamp 1666464484
transform 1 0 17756 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_189
timestamp 1666464484
transform 1 0 18492 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_193
timestamp 1666464484
transform 1 0 18860 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1666464484
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_197
timestamp 1666464484
transform 1 0 19228 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_205
timestamp 1666464484
transform 1 0 19964 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_213
timestamp 1666464484
transform 1 0 20700 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_221
timestamp 1666464484
transform 1 0 21436 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_229
timestamp 1666464484
transform 1 0 22172 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_237
timestamp 1666464484
transform 1 0 22908 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_245
timestamp 1666464484
transform 1 0 23644 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_249
timestamp 1666464484
transform 1 0 24012 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1666464484
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_253
timestamp 1666464484
transform 1 0 24380 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_261
timestamp 1666464484
transform 1 0 25116 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_269
timestamp 1666464484
transform 1 0 25852 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_277
timestamp 1666464484
transform 1 0 26588 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_285
timestamp 1666464484
transform 1 0 27324 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_293
timestamp 1666464484
transform 1 0 28060 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_301
timestamp 1666464484
transform 1 0 28796 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_305
timestamp 1666464484
transform 1 0 29164 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1666464484
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_309
timestamp 1666464484
transform 1 0 29532 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_317
timestamp 1666464484
transform 1 0 30268 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_325
timestamp 1666464484
transform 1 0 31004 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_333
timestamp 1666464484
transform 1 0 31740 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_341
timestamp 1666464484
transform 1 0 32476 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_349
timestamp 1666464484
transform 1 0 33212 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_357
timestamp 1666464484
transform 1 0 33948 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_362
timestamp 1666464484
transform 1 0 34408 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_90_365
timestamp 1666464484
transform 1 0 34684 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_373
timestamp 1666464484
transform 1 0 35420 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_381
timestamp 1666464484
transform 1 0 36156 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_389
timestamp 1666464484
transform 1 0 36892 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_397
timestamp 1666464484
transform 1 0 37628 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_405
timestamp 1666464484
transform 1 0 38364 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_413
timestamp 1666464484
transform 1 0 39100 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_417
timestamp 1666464484
transform 1 0 39468 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1666464484
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_421
timestamp 1666464484
transform 1 0 39836 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_429
timestamp 1666464484
transform 1 0 40572 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_437
timestamp 1666464484
transform 1 0 41308 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_445
timestamp 1666464484
transform 1 0 42044 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_453
timestamp 1666464484
transform 1 0 42780 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_461
timestamp 1666464484
transform 1 0 43516 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_469
timestamp 1666464484
transform 1 0 44252 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_473
timestamp 1666464484
transform 1 0 44620 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1666464484
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_477
timestamp 1666464484
transform 1 0 44988 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_485
timestamp 1666464484
transform 1 0 45724 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_493
timestamp 1666464484
transform 1 0 46460 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_501
timestamp 1666464484
transform 1 0 47196 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_509
timestamp 1666464484
transform 1 0 47932 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_517
timestamp 1666464484
transform 1 0 48668 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_525
timestamp 1666464484
transform 1 0 49404 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_529
timestamp 1666464484
transform 1 0 49772 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1666464484
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_533
timestamp 1666464484
transform 1 0 50140 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_541
timestamp 1666464484
transform 1 0 50876 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_549
timestamp 1666464484
transform 1 0 51612 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_557
timestamp 1666464484
transform 1 0 52348 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_565
timestamp 1666464484
transform 1 0 53084 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_573
timestamp 1666464484
transform 1 0 53820 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_581
timestamp 1666464484
transform 1 0 54556 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_585
timestamp 1666464484
transform 1 0 54924 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1666464484
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_90_589
timestamp 1666464484
transform 1 0 55292 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_597
timestamp 1666464484
transform 1 0 56028 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_605
timestamp 1666464484
transform 1 0 56764 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_90_613
timestamp 1666464484
transform 1 0 57500 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_90_621
timestamp 1666464484
transform 1 0 58236 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_91_3
timestamp 1666464484
transform 1 0 1380 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_11
timestamp 1666464484
transform 1 0 2116 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_19
timestamp 1666464484
transform 1 0 2852 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_27
timestamp 1666464484
transform 1 0 3588 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_35
timestamp 1666464484
transform 1 0 4324 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_43
timestamp 1666464484
transform 1 0 5060 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_51
timestamp 1666464484
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1666464484
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_57
timestamp 1666464484
transform 1 0 6348 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_65
timestamp 1666464484
transform 1 0 7084 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_73
timestamp 1666464484
transform 1 0 7820 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_81
timestamp 1666464484
transform 1 0 8556 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_89
timestamp 1666464484
transform 1 0 9292 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_97
timestamp 1666464484
transform 1 0 10028 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_105
timestamp 1666464484
transform 1 0 10764 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_109
timestamp 1666464484
transform 1 0 11132 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1666464484
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_113
timestamp 1666464484
transform 1 0 11500 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_121
timestamp 1666464484
transform 1 0 12236 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_129
timestamp 1666464484
transform 1 0 12972 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_137
timestamp 1666464484
transform 1 0 13708 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_145
timestamp 1666464484
transform 1 0 14444 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_153
timestamp 1666464484
transform 1 0 15180 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_161
timestamp 1666464484
transform 1 0 15916 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_165
timestamp 1666464484
transform 1 0 16284 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1666464484
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_169
timestamp 1666464484
transform 1 0 16652 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_177
timestamp 1666464484
transform 1 0 17388 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_185
timestamp 1666464484
transform 1 0 18124 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_193
timestamp 1666464484
transform 1 0 18860 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_201
timestamp 1666464484
transform 1 0 19596 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_209
timestamp 1666464484
transform 1 0 20332 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_217
timestamp 1666464484
transform 1 0 21068 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_221
timestamp 1666464484
transform 1 0 21436 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1666464484
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_225
timestamp 1666464484
transform 1 0 21804 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_233
timestamp 1666464484
transform 1 0 22540 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_241
timestamp 1666464484
transform 1 0 23276 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_249
timestamp 1666464484
transform 1 0 24012 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_257
timestamp 1666464484
transform 1 0 24748 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_265
timestamp 1666464484
transform 1 0 25484 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_273
timestamp 1666464484
transform 1 0 26220 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_277
timestamp 1666464484
transform 1 0 26588 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1666464484
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_281
timestamp 1666464484
transform 1 0 26956 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_289
timestamp 1666464484
transform 1 0 27692 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_297
timestamp 1666464484
transform 1 0 28428 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_305
timestamp 1666464484
transform 1 0 29164 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_313
timestamp 1666464484
transform 1 0 29900 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_321
timestamp 1666464484
transform 1 0 30636 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_329
timestamp 1666464484
transform 1 0 31372 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_333
timestamp 1666464484
transform 1 0 31740 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1666464484
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_337
timestamp 1666464484
transform 1 0 32108 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_345
timestamp 1666464484
transform 1 0 32844 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_353
timestamp 1666464484
transform 1 0 33580 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_357
timestamp 1666464484
transform 1 0 33948 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_91_380
timestamp 1666464484
transform 1 0 36064 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_388
timestamp 1666464484
transform 1 0 36800 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_91_393
timestamp 1666464484
transform 1 0 37260 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_401
timestamp 1666464484
transform 1 0 37996 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_409
timestamp 1666464484
transform 1 0 38732 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_417
timestamp 1666464484
transform 1 0 39468 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_425
timestamp 1666464484
transform 1 0 40204 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_433
timestamp 1666464484
transform 1 0 40940 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_441
timestamp 1666464484
transform 1 0 41676 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_445
timestamp 1666464484
transform 1 0 42044 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1666464484
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_449
timestamp 1666464484
transform 1 0 42412 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_457
timestamp 1666464484
transform 1 0 43148 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_465
timestamp 1666464484
transform 1 0 43884 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_473
timestamp 1666464484
transform 1 0 44620 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_481
timestamp 1666464484
transform 1 0 45356 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_489
timestamp 1666464484
transform 1 0 46092 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_497
timestamp 1666464484
transform 1 0 46828 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_501
timestamp 1666464484
transform 1 0 47196 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1666464484
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_505
timestamp 1666464484
transform 1 0 47564 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_513
timestamp 1666464484
transform 1 0 48300 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_521
timestamp 1666464484
transform 1 0 49036 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_529
timestamp 1666464484
transform 1 0 49772 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_537
timestamp 1666464484
transform 1 0 50508 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_545
timestamp 1666464484
transform 1 0 51244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_553
timestamp 1666464484
transform 1 0 51980 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_557
timestamp 1666464484
transform 1 0 52348 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1666464484
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_561
timestamp 1666464484
transform 1 0 52716 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_569
timestamp 1666464484
transform 1 0 53452 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_577
timestamp 1666464484
transform 1 0 54188 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_585
timestamp 1666464484
transform 1 0 54924 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_593
timestamp 1666464484
transform 1 0 55660 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_91_601
timestamp 1666464484
transform 1 0 56396 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_91_609
timestamp 1666464484
transform 1 0 57132 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_613
timestamp 1666464484
transform 1 0 57500 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1666464484
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_91_617
timestamp 1666464484
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_3
timestamp 1666464484
transform 1 0 1380 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_11
timestamp 1666464484
transform 1 0 2116 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_19
timestamp 1666464484
transform 1 0 2852 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1666464484
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_29
timestamp 1666464484
transform 1 0 3772 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_37
timestamp 1666464484
transform 1 0 4508 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_45
timestamp 1666464484
transform 1 0 5244 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_53
timestamp 1666464484
transform 1 0 5980 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_61
timestamp 1666464484
transform 1 0 6716 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_69
timestamp 1666464484
transform 1 0 7452 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_77
timestamp 1666464484
transform 1 0 8188 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_81
timestamp 1666464484
transform 1 0 8556 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1666464484
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_85
timestamp 1666464484
transform 1 0 8924 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_93
timestamp 1666464484
transform 1 0 9660 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_101
timestamp 1666464484
transform 1 0 10396 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_109
timestamp 1666464484
transform 1 0 11132 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_117
timestamp 1666464484
transform 1 0 11868 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_125
timestamp 1666464484
transform 1 0 12604 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_133
timestamp 1666464484
transform 1 0 13340 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_137
timestamp 1666464484
transform 1 0 13708 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1666464484
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_141
timestamp 1666464484
transform 1 0 14076 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_149
timestamp 1666464484
transform 1 0 14812 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_157
timestamp 1666464484
transform 1 0 15548 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_165
timestamp 1666464484
transform 1 0 16284 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_173
timestamp 1666464484
transform 1 0 17020 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_181
timestamp 1666464484
transform 1 0 17756 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_189
timestamp 1666464484
transform 1 0 18492 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_193
timestamp 1666464484
transform 1 0 18860 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1666464484
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_197
timestamp 1666464484
transform 1 0 19228 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_205
timestamp 1666464484
transform 1 0 19964 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_213
timestamp 1666464484
transform 1 0 20700 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_221
timestamp 1666464484
transform 1 0 21436 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_229
timestamp 1666464484
transform 1 0 22172 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_237
timestamp 1666464484
transform 1 0 22908 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_245
timestamp 1666464484
transform 1 0 23644 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_249
timestamp 1666464484
transform 1 0 24012 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1666464484
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_253
timestamp 1666464484
transform 1 0 24380 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_261
timestamp 1666464484
transform 1 0 25116 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_269
timestamp 1666464484
transform 1 0 25852 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_277
timestamp 1666464484
transform 1 0 26588 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_285
timestamp 1666464484
transform 1 0 27324 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_293
timestamp 1666464484
transform 1 0 28060 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_301
timestamp 1666464484
transform 1 0 28796 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_305
timestamp 1666464484
transform 1 0 29164 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1666464484
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_309
timestamp 1666464484
transform 1 0 29532 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_317
timestamp 1666464484
transform 1 0 30268 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_325
timestamp 1666464484
transform 1 0 31004 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_333
timestamp 1666464484
transform 1 0 31740 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_92_339
timestamp 1666464484
transform 1 0 32292 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_347
timestamp 1666464484
transform 1 0 33028 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_355
timestamp 1666464484
transform 1 0 33764 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1666464484
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_365
timestamp 1666464484
transform 1 0 34684 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_373
timestamp 1666464484
transform 1 0 35420 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_381
timestamp 1666464484
transform 1 0 36156 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_389
timestamp 1666464484
transform 1 0 36892 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_397
timestamp 1666464484
transform 1 0 37628 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_405
timestamp 1666464484
transform 1 0 38364 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_413
timestamp 1666464484
transform 1 0 39100 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_417
timestamp 1666464484
transform 1 0 39468 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1666464484
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_421
timestamp 1666464484
transform 1 0 39836 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_429
timestamp 1666464484
transform 1 0 40572 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_437
timestamp 1666464484
transform 1 0 41308 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_445
timestamp 1666464484
transform 1 0 42044 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_453
timestamp 1666464484
transform 1 0 42780 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_461
timestamp 1666464484
transform 1 0 43516 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_469
timestamp 1666464484
transform 1 0 44252 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_473
timestamp 1666464484
transform 1 0 44620 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1666464484
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_477
timestamp 1666464484
transform 1 0 44988 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_485
timestamp 1666464484
transform 1 0 45724 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_493
timestamp 1666464484
transform 1 0 46460 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_501
timestamp 1666464484
transform 1 0 47196 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_509
timestamp 1666464484
transform 1 0 47932 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_517
timestamp 1666464484
transform 1 0 48668 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_525
timestamp 1666464484
transform 1 0 49404 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_529
timestamp 1666464484
transform 1 0 49772 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1666464484
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_533
timestamp 1666464484
transform 1 0 50140 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_541
timestamp 1666464484
transform 1 0 50876 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_549
timestamp 1666464484
transform 1 0 51612 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_557
timestamp 1666464484
transform 1 0 52348 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_565
timestamp 1666464484
transform 1 0 53084 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_573
timestamp 1666464484
transform 1 0 53820 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_581
timestamp 1666464484
transform 1 0 54556 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_585
timestamp 1666464484
transform 1 0 54924 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1666464484
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_92_589
timestamp 1666464484
transform 1 0 55292 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_597
timestamp 1666464484
transform 1 0 56028 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_605
timestamp 1666464484
transform 1 0 56764 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_92_613
timestamp 1666464484
transform 1 0 57500 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_92_621
timestamp 1666464484
transform 1 0 58236 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_93_3
timestamp 1666464484
transform 1 0 1380 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_11
timestamp 1666464484
transform 1 0 2116 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_19
timestamp 1666464484
transform 1 0 2852 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_27
timestamp 1666464484
transform 1 0 3588 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_35
timestamp 1666464484
transform 1 0 4324 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_43
timestamp 1666464484
transform 1 0 5060 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_51
timestamp 1666464484
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1666464484
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_57
timestamp 1666464484
transform 1 0 6348 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_65
timestamp 1666464484
transform 1 0 7084 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_73
timestamp 1666464484
transform 1 0 7820 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_81
timestamp 1666464484
transform 1 0 8556 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_89
timestamp 1666464484
transform 1 0 9292 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_97
timestamp 1666464484
transform 1 0 10028 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_105
timestamp 1666464484
transform 1 0 10764 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_109
timestamp 1666464484
transform 1 0 11132 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1666464484
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_113
timestamp 1666464484
transform 1 0 11500 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_121
timestamp 1666464484
transform 1 0 12236 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_129
timestamp 1666464484
transform 1 0 12972 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_137
timestamp 1666464484
transform 1 0 13708 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_145
timestamp 1666464484
transform 1 0 14444 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_153
timestamp 1666464484
transform 1 0 15180 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_161
timestamp 1666464484
transform 1 0 15916 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_165
timestamp 1666464484
transform 1 0 16284 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1666464484
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_169
timestamp 1666464484
transform 1 0 16652 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_177
timestamp 1666464484
transform 1 0 17388 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_185
timestamp 1666464484
transform 1 0 18124 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_193
timestamp 1666464484
transform 1 0 18860 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_201
timestamp 1666464484
transform 1 0 19596 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_209
timestamp 1666464484
transform 1 0 20332 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_217
timestamp 1666464484
transform 1 0 21068 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_221
timestamp 1666464484
transform 1 0 21436 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1666464484
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_225
timestamp 1666464484
transform 1 0 21804 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_233
timestamp 1666464484
transform 1 0 22540 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_241
timestamp 1666464484
transform 1 0 23276 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_249
timestamp 1666464484
transform 1 0 24012 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_257
timestamp 1666464484
transform 1 0 24748 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_265
timestamp 1666464484
transform 1 0 25484 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_273
timestamp 1666464484
transform 1 0 26220 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_277
timestamp 1666464484
transform 1 0 26588 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1666464484
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_281
timestamp 1666464484
transform 1 0 26956 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_289
timestamp 1666464484
transform 1 0 27692 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_297
timestamp 1666464484
transform 1 0 28428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_305
timestamp 1666464484
transform 1 0 29164 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_313
timestamp 1666464484
transform 1 0 29900 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_317
timestamp 1666464484
transform 1 0 30268 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_93_321
timestamp 1666464484
transform 1 0 30636 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_329
timestamp 1666464484
transform 1 0 31372 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_93_332
timestamp 1666464484
transform 1 0 31648 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_93_337
timestamp 1666464484
transform 1 0 32108 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_341
timestamp 1666464484
transform 1 0 32476 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_343
timestamp 1666464484
transform 1 0 32660 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_93_346
timestamp 1666464484
transform 1 0 32936 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_93_352
timestamp 1666464484
transform 1 0 33488 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_93_358
timestamp 1666464484
transform 1 0 34040 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_93_364
timestamp 1666464484
transform 1 0 34592 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_372
timestamp 1666464484
transform 1 0 35328 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_380
timestamp 1666464484
transform 1 0 36064 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_388
timestamp 1666464484
transform 1 0 36800 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_93_393
timestamp 1666464484
transform 1 0 37260 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_401
timestamp 1666464484
transform 1 0 37996 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_409
timestamp 1666464484
transform 1 0 38732 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_417
timestamp 1666464484
transform 1 0 39468 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_93_423
timestamp 1666464484
transform 1 0 40020 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_431
timestamp 1666464484
transform 1 0 40756 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_439
timestamp 1666464484
transform 1 0 41492 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1666464484
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_449
timestamp 1666464484
transform 1 0 42412 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_457
timestamp 1666464484
transform 1 0 43148 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_465
timestamp 1666464484
transform 1 0 43884 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_473
timestamp 1666464484
transform 1 0 44620 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_481
timestamp 1666464484
transform 1 0 45356 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_489
timestamp 1666464484
transform 1 0 46092 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_497
timestamp 1666464484
transform 1 0 46828 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_501
timestamp 1666464484
transform 1 0 47196 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1666464484
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_505
timestamp 1666464484
transform 1 0 47564 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_513
timestamp 1666464484
transform 1 0 48300 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_521
timestamp 1666464484
transform 1 0 49036 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_529
timestamp 1666464484
transform 1 0 49772 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_537
timestamp 1666464484
transform 1 0 50508 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_545
timestamp 1666464484
transform 1 0 51244 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_553
timestamp 1666464484
transform 1 0 51980 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_557
timestamp 1666464484
transform 1 0 52348 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1666464484
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_561
timestamp 1666464484
transform 1 0 52716 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_569
timestamp 1666464484
transform 1 0 53452 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_577
timestamp 1666464484
transform 1 0 54188 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_585
timestamp 1666464484
transform 1 0 54924 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_593
timestamp 1666464484
transform 1 0 55660 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_93_601
timestamp 1666464484
transform 1 0 56396 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_93_609
timestamp 1666464484
transform 1 0 57132 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_613
timestamp 1666464484
transform 1 0 57500 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1666464484
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_93_617
timestamp 1666464484
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_3
timestamp 1666464484
transform 1 0 1380 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_11
timestamp 1666464484
transform 1 0 2116 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_19
timestamp 1666464484
transform 1 0 2852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1666464484
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_29
timestamp 1666464484
transform 1 0 3772 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_37
timestamp 1666464484
transform 1 0 4508 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_45
timestamp 1666464484
transform 1 0 5244 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_53
timestamp 1666464484
transform 1 0 5980 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_61
timestamp 1666464484
transform 1 0 6716 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_69
timestamp 1666464484
transform 1 0 7452 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_77
timestamp 1666464484
transform 1 0 8188 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_81
timestamp 1666464484
transform 1 0 8556 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1666464484
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_85
timestamp 1666464484
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_93
timestamp 1666464484
transform 1 0 9660 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_101
timestamp 1666464484
transform 1 0 10396 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_109
timestamp 1666464484
transform 1 0 11132 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_117
timestamp 1666464484
transform 1 0 11868 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_125
timestamp 1666464484
transform 1 0 12604 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_133
timestamp 1666464484
transform 1 0 13340 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_137
timestamp 1666464484
transform 1 0 13708 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1666464484
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_141
timestamp 1666464484
transform 1 0 14076 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_149
timestamp 1666464484
transform 1 0 14812 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_157
timestamp 1666464484
transform 1 0 15548 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_165
timestamp 1666464484
transform 1 0 16284 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_173
timestamp 1666464484
transform 1 0 17020 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_181
timestamp 1666464484
transform 1 0 17756 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_189
timestamp 1666464484
transform 1 0 18492 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_193
timestamp 1666464484
transform 1 0 18860 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1666464484
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_197
timestamp 1666464484
transform 1 0 19228 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_205
timestamp 1666464484
transform 1 0 19964 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_213
timestamp 1666464484
transform 1 0 20700 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_221
timestamp 1666464484
transform 1 0 21436 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_229
timestamp 1666464484
transform 1 0 22172 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_237
timestamp 1666464484
transform 1 0 22908 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_245
timestamp 1666464484
transform 1 0 23644 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_249
timestamp 1666464484
transform 1 0 24012 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1666464484
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_253
timestamp 1666464484
transform 1 0 24380 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_261
timestamp 1666464484
transform 1 0 25116 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_269
timestamp 1666464484
transform 1 0 25852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_277
timestamp 1666464484
transform 1 0 26588 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_279
timestamp 1666464484
transform 1 0 26772 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_282
timestamp 1666464484
transform 1 0 27048 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_290
timestamp 1666464484
transform 1 0 27784 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_293
timestamp 1666464484
transform 1 0 28060 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_301
timestamp 1666464484
transform 1 0 28796 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_303
timestamp 1666464484
transform 1 0 28980 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_306
timestamp 1666464484
transform 1 0 29256 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_94_309
timestamp 1666464484
transform 1 0 29532 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_94_318
timestamp 1666464484
transform 1 0 30360 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_94_324
timestamp 1666464484
transform 1 0 30912 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_328
timestamp 1666464484
transform 1 0 31280 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_94_331
timestamp 1666464484
transform 1 0 31556 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_94_341
timestamp 1666464484
transform 1 0 32476 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_94_351
timestamp 1666464484
transform 1 0 33396 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_355
timestamp 1666464484
transform 1 0 33764 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_362
timestamp 1666464484
transform 1 0 34408 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_365
timestamp 1666464484
transform 1 0 34684 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_94_373
timestamp 1666464484
transform 1 0 35420 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_94_379
timestamp 1666464484
transform 1 0 35972 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_387
timestamp 1666464484
transform 1 0 36708 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_395
timestamp 1666464484
transform 1 0 37444 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_403
timestamp 1666464484
transform 1 0 38180 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_411
timestamp 1666464484
transform 1 0 38916 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_417
timestamp 1666464484
transform 1 0 39468 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1666464484
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_421
timestamp 1666464484
transform 1 0 39836 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_423
timestamp 1666464484
transform 1 0 40020 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_94_426
timestamp 1666464484
transform 1 0 40296 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_430
timestamp 1666464484
transform 1 0 40664 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_94_433
timestamp 1666464484
transform 1 0 40940 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_94_439
timestamp 1666464484
transform 1 0 41492 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_443
timestamp 1666464484
transform 1 0 41860 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_94_450
timestamp 1666464484
transform 1 0 42504 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_458
timestamp 1666464484
transform 1 0 43240 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_466
timestamp 1666464484
transform 1 0 43976 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_474
timestamp 1666464484
transform 1 0 44712 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_94_477
timestamp 1666464484
transform 1 0 44988 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_485
timestamp 1666464484
transform 1 0 45724 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_493
timestamp 1666464484
transform 1 0 46460 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_501
timestamp 1666464484
transform 1 0 47196 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_509
timestamp 1666464484
transform 1 0 47932 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_517
timestamp 1666464484
transform 1 0 48668 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_525
timestamp 1666464484
transform 1 0 49404 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_529
timestamp 1666464484
transform 1 0 49772 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1666464484
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_533
timestamp 1666464484
transform 1 0 50140 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_541
timestamp 1666464484
transform 1 0 50876 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_549
timestamp 1666464484
transform 1 0 51612 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_557
timestamp 1666464484
transform 1 0 52348 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_565
timestamp 1666464484
transform 1 0 53084 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_573
timestamp 1666464484
transform 1 0 53820 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_581
timestamp 1666464484
transform 1 0 54556 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_585
timestamp 1666464484
transform 1 0 54924 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1666464484
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_94_589
timestamp 1666464484
transform 1 0 55292 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_597
timestamp 1666464484
transform 1 0 56028 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_605
timestamp 1666464484
transform 1 0 56764 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_94_613
timestamp 1666464484
transform 1 0 57500 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_94_621
timestamp 1666464484
transform 1 0 58236 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_95_3
timestamp 1666464484
transform 1 0 1380 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_11
timestamp 1666464484
transform 1 0 2116 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_19
timestamp 1666464484
transform 1 0 2852 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_27
timestamp 1666464484
transform 1 0 3588 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_35
timestamp 1666464484
transform 1 0 4324 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_43
timestamp 1666464484
transform 1 0 5060 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_51
timestamp 1666464484
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1666464484
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_95_57
timestamp 1666464484
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_65
timestamp 1666464484
transform 1 0 7084 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_73
timestamp 1666464484
transform 1 0 7820 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_81
timestamp 1666464484
transform 1 0 8556 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_89
timestamp 1666464484
transform 1 0 9292 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_97
timestamp 1666464484
transform 1 0 10028 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_105
timestamp 1666464484
transform 1 0 10764 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_109
timestamp 1666464484
transform 1 0 11132 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1666464484
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_95_113
timestamp 1666464484
transform 1 0 11500 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_121
timestamp 1666464484
transform 1 0 12236 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_129
timestamp 1666464484
transform 1 0 12972 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_137
timestamp 1666464484
transform 1 0 13708 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_145
timestamp 1666464484
transform 1 0 14444 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_153
timestamp 1666464484
transform 1 0 15180 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_161
timestamp 1666464484
transform 1 0 15916 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_165
timestamp 1666464484
transform 1 0 16284 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1666464484
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_95_169
timestamp 1666464484
transform 1 0 16652 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_177
timestamp 1666464484
transform 1 0 17388 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_185
timestamp 1666464484
transform 1 0 18124 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_193
timestamp 1666464484
transform 1 0 18860 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_201
timestamp 1666464484
transform 1 0 19596 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_209
timestamp 1666464484
transform 1 0 20332 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_217
timestamp 1666464484
transform 1 0 21068 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_221
timestamp 1666464484
transform 1 0 21436 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1666464484
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_95_225
timestamp 1666464484
transform 1 0 21804 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_233
timestamp 1666464484
transform 1 0 22540 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_241
timestamp 1666464484
transform 1 0 23276 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_249
timestamp 1666464484
transform 1 0 24012 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_257
timestamp 1666464484
transform 1 0 24748 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_265
timestamp 1666464484
transform 1 0 25484 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_273
timestamp 1666464484
transform 1 0 26220 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_275
timestamp 1666464484
transform 1 0 26404 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_278
timestamp 1666464484
transform 1 0 26680 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_281
timestamp 1666464484
transform 1 0 26956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_95_285
timestamp 1666464484
transform 1 0 27324 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_291
timestamp 1666464484
transform 1 0 27876 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_302
timestamp 1666464484
transform 1 0 28888 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_306
timestamp 1666464484
transform 1 0 29256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_95_312
timestamp 1666464484
transform 1 0 29808 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_323
timestamp 1666464484
transform 1 0 30820 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_329
timestamp 1666464484
transform 1 0 31372 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_333
timestamp 1666464484
transform 1 0 31740 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1666464484
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_337
timestamp 1666464484
transform 1 0 32108 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_95_346
timestamp 1666464484
transform 1 0 32936 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_362
timestamp 1666464484
transform 1 0 34408 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_373
timestamp 1666464484
transform 1 0 35420 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_379
timestamp 1666464484
transform 1 0 35972 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_385
timestamp 1666464484
transform 1 0 36524 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_389
timestamp 1666464484
transform 1 0 36892 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1666464484
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_393
timestamp 1666464484
transform 1 0 37260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_95_397
timestamp 1666464484
transform 1 0 37628 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_405
timestamp 1666464484
transform 1 0 38364 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_409
timestamp 1666464484
transform 1 0 38732 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_411
timestamp 1666464484
transform 1 0 38916 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_95_415
timestamp 1666464484
transform 1 0 39284 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_422
timestamp 1666464484
transform 1 0 39928 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_429
timestamp 1666464484
transform 1 0 40572 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_95_440
timestamp 1666464484
transform 1 0 41584 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_446
timestamp 1666464484
transform 1 0 42136 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_449
timestamp 1666464484
transform 1 0 42412 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_95_457
timestamp 1666464484
transform 1 0 43148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_461
timestamp 1666464484
transform 1 0 43516 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_95_469
timestamp 1666464484
transform 1 0 44252 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_477
timestamp 1666464484
transform 1 0 44988 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_485
timestamp 1666464484
transform 1 0 45724 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_493
timestamp 1666464484
transform 1 0 46460 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_501
timestamp 1666464484
transform 1 0 47196 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1666464484
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_95_505
timestamp 1666464484
transform 1 0 47564 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_513
timestamp 1666464484
transform 1 0 48300 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_521
timestamp 1666464484
transform 1 0 49036 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_529
timestamp 1666464484
transform 1 0 49772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_537
timestamp 1666464484
transform 1 0 50508 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_545
timestamp 1666464484
transform 1 0 51244 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_553
timestamp 1666464484
transform 1 0 51980 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_557
timestamp 1666464484
transform 1 0 52348 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1666464484
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_95_561
timestamp 1666464484
transform 1 0 52716 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_569
timestamp 1666464484
transform 1 0 53452 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_577
timestamp 1666464484
transform 1 0 54188 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_585
timestamp 1666464484
transform 1 0 54924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_593
timestamp 1666464484
transform 1 0 55660 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_95_601
timestamp 1666464484
transform 1 0 56396 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_95_609
timestamp 1666464484
transform 1 0 57132 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_613
timestamp 1666464484
transform 1 0 57500 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1666464484
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_95_617
timestamp 1666464484
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_3
timestamp 1666464484
transform 1 0 1380 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_11
timestamp 1666464484
transform 1 0 2116 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_19
timestamp 1666464484
transform 1 0 2852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1666464484
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_96_29
timestamp 1666464484
transform 1 0 3772 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_37
timestamp 1666464484
transform 1 0 4508 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_45
timestamp 1666464484
transform 1 0 5244 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_53
timestamp 1666464484
transform 1 0 5980 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_61
timestamp 1666464484
transform 1 0 6716 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_69
timestamp 1666464484
transform 1 0 7452 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_77
timestamp 1666464484
transform 1 0 8188 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_81
timestamp 1666464484
transform 1 0 8556 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1666464484
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_96_85
timestamp 1666464484
transform 1 0 8924 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_93
timestamp 1666464484
transform 1 0 9660 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_101
timestamp 1666464484
transform 1 0 10396 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_109
timestamp 1666464484
transform 1 0 11132 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_117
timestamp 1666464484
transform 1 0 11868 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_125
timestamp 1666464484
transform 1 0 12604 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_133
timestamp 1666464484
transform 1 0 13340 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_137
timestamp 1666464484
transform 1 0 13708 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1666464484
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_96_141
timestamp 1666464484
transform 1 0 14076 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_149
timestamp 1666464484
transform 1 0 14812 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_157
timestamp 1666464484
transform 1 0 15548 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_165
timestamp 1666464484
transform 1 0 16284 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_173
timestamp 1666464484
transform 1 0 17020 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_181
timestamp 1666464484
transform 1 0 17756 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_189
timestamp 1666464484
transform 1 0 18492 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_193
timestamp 1666464484
transform 1 0 18860 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1666464484
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_96_197
timestamp 1666464484
transform 1 0 19228 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_205
timestamp 1666464484
transform 1 0 19964 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_213
timestamp 1666464484
transform 1 0 20700 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_221
timestamp 1666464484
transform 1 0 21436 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_229
timestamp 1666464484
transform 1 0 22172 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_237
timestamp 1666464484
transform 1 0 22908 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_245
timestamp 1666464484
transform 1 0 23644 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_249
timestamp 1666464484
transform 1 0 24012 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1666464484
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_96_253
timestamp 1666464484
transform 1 0 24380 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_257
timestamp 1666464484
transform 1 0 24748 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_259
timestamp 1666464484
transform 1 0 24932 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_96_262
timestamp 1666464484
transform 1 0 25208 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_266
timestamp 1666464484
transform 1 0 25576 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_96_270
timestamp 1666464484
transform 1 0 25944 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_277
timestamp 1666464484
transform 1 0 26588 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_284
timestamp 1666464484
transform 1 0 27232 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_288
timestamp 1666464484
transform 1 0 27600 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_96_292
timestamp 1666464484
transform 1 0 27968 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_302
timestamp 1666464484
transform 1 0 28888 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_306
timestamp 1666464484
transform 1 0 29256 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_309
timestamp 1666464484
transform 1 0 29532 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_96_318
timestamp 1666464484
transform 1 0 30360 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_322
timestamp 1666464484
transform 1 0 30728 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_96_327
timestamp 1666464484
transform 1 0 31188 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_331
timestamp 1666464484
transform 1 0 31556 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_96_339
timestamp 1666464484
transform 1 0 32292 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_349
timestamp 1666464484
transform 1 0 33212 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_358
timestamp 1666464484
transform 1 0 34040 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_362
timestamp 1666464484
transform 1 0 34408 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_365
timestamp 1666464484
transform 1 0 34684 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_96_370
timestamp 1666464484
transform 1 0 35144 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_376
timestamp 1666464484
transform 1 0 35696 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_382
timestamp 1666464484
transform 1 0 36248 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_388
timestamp 1666464484
transform 1 0 36800 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_96_394
timestamp 1666464484
transform 1 0 37352 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_407
timestamp 1666464484
transform 1 0 38548 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_418
timestamp 1666464484
transform 1 0 39560 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_421
timestamp 1666464484
transform 1 0 39836 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_96_426
timestamp 1666464484
transform 1 0 40296 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_430
timestamp 1666464484
transform 1 0 40664 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_96_437
timestamp 1666464484
transform 1 0 41308 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_447
timestamp 1666464484
transform 1 0 42228 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_459
timestamp 1666464484
transform 1 0 43332 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_96_470
timestamp 1666464484
transform 1 0 44344 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_474
timestamp 1666464484
transform 1 0 44712 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_96_477
timestamp 1666464484
transform 1 0 44988 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_485
timestamp 1666464484
transform 1 0 45724 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_493
timestamp 1666464484
transform 1 0 46460 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_501
timestamp 1666464484
transform 1 0 47196 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_509
timestamp 1666464484
transform 1 0 47932 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_517
timestamp 1666464484
transform 1 0 48668 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_525
timestamp 1666464484
transform 1 0 49404 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_529
timestamp 1666464484
transform 1 0 49772 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1666464484
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_96_533
timestamp 1666464484
transform 1 0 50140 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_541
timestamp 1666464484
transform 1 0 50876 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_549
timestamp 1666464484
transform 1 0 51612 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_557
timestamp 1666464484
transform 1 0 52348 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_565
timestamp 1666464484
transform 1 0 53084 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_573
timestamp 1666464484
transform 1 0 53820 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_581
timestamp 1666464484
transform 1 0 54556 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_585
timestamp 1666464484
transform 1 0 54924 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1666464484
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_96_589
timestamp 1666464484
transform 1 0 55292 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_597
timestamp 1666464484
transform 1 0 56028 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_605
timestamp 1666464484
transform 1 0 56764 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_96_613
timestamp 1666464484
transform 1 0 57500 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_96_621
timestamp 1666464484
transform 1 0 58236 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_97_3
timestamp 1666464484
transform 1 0 1380 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_11
timestamp 1666464484
transform 1 0 2116 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_19
timestamp 1666464484
transform 1 0 2852 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_27
timestamp 1666464484
transform 1 0 3588 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_35
timestamp 1666464484
transform 1 0 4324 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_43
timestamp 1666464484
transform 1 0 5060 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_51
timestamp 1666464484
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1666464484
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_97_57
timestamp 1666464484
transform 1 0 6348 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_65
timestamp 1666464484
transform 1 0 7084 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_73
timestamp 1666464484
transform 1 0 7820 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_81
timestamp 1666464484
transform 1 0 8556 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_89
timestamp 1666464484
transform 1 0 9292 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_97
timestamp 1666464484
transform 1 0 10028 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_105
timestamp 1666464484
transform 1 0 10764 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_109
timestamp 1666464484
transform 1 0 11132 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1666464484
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_97_113
timestamp 1666464484
transform 1 0 11500 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_121
timestamp 1666464484
transform 1 0 12236 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_129
timestamp 1666464484
transform 1 0 12972 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_137
timestamp 1666464484
transform 1 0 13708 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_145
timestamp 1666464484
transform 1 0 14444 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_153
timestamp 1666464484
transform 1 0 15180 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_161
timestamp 1666464484
transform 1 0 15916 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_165
timestamp 1666464484
transform 1 0 16284 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1666464484
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_97_169
timestamp 1666464484
transform 1 0 16652 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_177
timestamp 1666464484
transform 1 0 17388 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_185
timestamp 1666464484
transform 1 0 18124 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_193
timestamp 1666464484
transform 1 0 18860 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_201
timestamp 1666464484
transform 1 0 19596 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_209
timestamp 1666464484
transform 1 0 20332 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_217
timestamp 1666464484
transform 1 0 21068 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_221
timestamp 1666464484
transform 1 0 21436 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1666464484
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_97_225
timestamp 1666464484
transform 1 0 21804 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_233
timestamp 1666464484
transform 1 0 22540 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_241
timestamp 1666464484
transform 1 0 23276 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_245
timestamp 1666464484
transform 1 0 23644 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_97_249
timestamp 1666464484
transform 1 0 24012 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_255
timestamp 1666464484
transform 1 0 24564 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_261
timestamp 1666464484
transform 1 0 25116 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_268
timestamp 1666464484
transform 1 0 25760 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_272
timestamp 1666464484
transform 1 0 26128 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_274
timestamp 1666464484
transform 1 0 26312 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_278
timestamp 1666464484
transform 1 0 26680 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_281
timestamp 1666464484
transform 1 0 26956 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_97_286
timestamp 1666464484
transform 1 0 27416 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_293
timestamp 1666464484
transform 1 0 28060 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_300
timestamp 1666464484
transform 1 0 28704 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_308
timestamp 1666464484
transform 1 0 29440 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_317
timestamp 1666464484
transform 1 0 30268 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_321
timestamp 1666464484
transform 1 0 30636 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_323
timestamp 1666464484
transform 1 0 30820 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_97_329
timestamp 1666464484
transform 1 0 31372 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_333
timestamp 1666464484
transform 1 0 31740 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1666464484
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_337
timestamp 1666464484
transform 1 0 32108 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_97_344
timestamp 1666464484
transform 1 0 32752 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_351
timestamp 1666464484
transform 1 0 33396 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_358
timestamp 1666464484
transform 1 0 34040 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_365
timestamp 1666464484
transform 1 0 34684 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_376
timestamp 1666464484
transform 1 0 35696 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_383
timestamp 1666464484
transform 1 0 36340 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_390
timestamp 1666464484
transform 1 0 36984 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_393
timestamp 1666464484
transform 1 0 37260 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_97_398
timestamp 1666464484
transform 1 0 37720 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_402
timestamp 1666464484
transform 1 0 38088 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_97_410
timestamp 1666464484
transform 1 0 38824 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_419
timestamp 1666464484
transform 1 0 39652 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_427
timestamp 1666464484
transform 1 0 40388 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_433
timestamp 1666464484
transform 1 0 40940 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_443
timestamp 1666464484
transform 1 0 41860 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1666464484
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_449
timestamp 1666464484
transform 1 0 42412 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_451
timestamp 1666464484
transform 1 0 42596 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_97_458
timestamp 1666464484
transform 1 0 43240 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_465
timestamp 1666464484
transform 1 0 43884 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_472
timestamp 1666464484
transform 1 0 44528 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_97_478
timestamp 1666464484
transform 1 0 45080 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_482
timestamp 1666464484
transform 1 0 45448 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_97_486
timestamp 1666464484
transform 1 0 45816 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_97_492
timestamp 1666464484
transform 1 0 46368 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_500
timestamp 1666464484
transform 1 0 47104 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_97_505
timestamp 1666464484
transform 1 0 47564 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_513
timestamp 1666464484
transform 1 0 48300 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_521
timestamp 1666464484
transform 1 0 49036 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_529
timestamp 1666464484
transform 1 0 49772 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_537
timestamp 1666464484
transform 1 0 50508 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_545
timestamp 1666464484
transform 1 0 51244 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_553
timestamp 1666464484
transform 1 0 51980 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_557
timestamp 1666464484
transform 1 0 52348 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1666464484
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_97_561
timestamp 1666464484
transform 1 0 52716 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_569
timestamp 1666464484
transform 1 0 53452 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_577
timestamp 1666464484
transform 1 0 54188 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_585
timestamp 1666464484
transform 1 0 54924 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_593
timestamp 1666464484
transform 1 0 55660 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_97_601
timestamp 1666464484
transform 1 0 56396 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_97_609
timestamp 1666464484
transform 1 0 57132 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_613
timestamp 1666464484
transform 1 0 57500 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1666464484
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_97_617
timestamp 1666464484
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_3
timestamp 1666464484
transform 1 0 1380 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_11
timestamp 1666464484
transform 1 0 2116 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_19
timestamp 1666464484
transform 1 0 2852 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1666464484
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_98_29
timestamp 1666464484
transform 1 0 3772 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_37
timestamp 1666464484
transform 1 0 4508 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_45
timestamp 1666464484
transform 1 0 5244 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_53
timestamp 1666464484
transform 1 0 5980 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_61
timestamp 1666464484
transform 1 0 6716 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_69
timestamp 1666464484
transform 1 0 7452 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_98_77
timestamp 1666464484
transform 1 0 8188 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_81
timestamp 1666464484
transform 1 0 8556 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1666464484
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_98_85
timestamp 1666464484
transform 1 0 8924 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_93
timestamp 1666464484
transform 1 0 9660 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_101
timestamp 1666464484
transform 1 0 10396 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_109
timestamp 1666464484
transform 1 0 11132 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_117
timestamp 1666464484
transform 1 0 11868 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_125
timestamp 1666464484
transform 1 0 12604 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_98_133
timestamp 1666464484
transform 1 0 13340 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_137
timestamp 1666464484
transform 1 0 13708 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1666464484
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_98_141
timestamp 1666464484
transform 1 0 14076 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_149
timestamp 1666464484
transform 1 0 14812 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_157
timestamp 1666464484
transform 1 0 15548 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_165
timestamp 1666464484
transform 1 0 16284 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_173
timestamp 1666464484
transform 1 0 17020 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_181
timestamp 1666464484
transform 1 0 17756 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_98_189
timestamp 1666464484
transform 1 0 18492 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_193
timestamp 1666464484
transform 1 0 18860 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1666464484
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_98_197
timestamp 1666464484
transform 1 0 19228 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_205
timestamp 1666464484
transform 1 0 19964 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_213
timestamp 1666464484
transform 1 0 20700 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_221
timestamp 1666464484
transform 1 0 21436 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_229
timestamp 1666464484
transform 1 0 22172 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_98_237
timestamp 1666464484
transform 1 0 22908 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_243
timestamp 1666464484
transform 1 0 23460 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_250
timestamp 1666464484
transform 1 0 24104 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_253
timestamp 1666464484
transform 1 0 24380 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_255
timestamp 1666464484
transform 1 0 24564 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_98_259
timestamp 1666464484
transform 1 0 24932 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_268
timestamp 1666464484
transform 1 0 25760 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_274
timestamp 1666464484
transform 1 0 26312 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_283
timestamp 1666464484
transform 1 0 27140 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_287
timestamp 1666464484
transform 1 0 27508 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_98_293
timestamp 1666464484
transform 1 0 28060 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_304
timestamp 1666464484
transform 1 0 29072 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_309
timestamp 1666464484
transform 1 0 29532 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_318
timestamp 1666464484
transform 1 0 30360 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_322
timestamp 1666464484
transform 1 0 30728 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_98_332
timestamp 1666464484
transform 1 0 31648 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_342
timestamp 1666464484
transform 1 0 32568 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_352
timestamp 1666464484
transform 1 0 33488 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_356
timestamp 1666464484
transform 1 0 33856 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_362
timestamp 1666464484
transform 1 0 34408 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_365
timestamp 1666464484
transform 1 0 34684 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_98_374
timestamp 1666464484
transform 1 0 35512 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_381
timestamp 1666464484
transform 1 0 36156 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_392
timestamp 1666464484
transform 1 0 37168 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_398
timestamp 1666464484
transform 1 0 37720 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_408
timestamp 1666464484
transform 1 0 38640 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_417
timestamp 1666464484
transform 1 0 39468 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1666464484
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_421
timestamp 1666464484
transform 1 0 39836 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_98_428
timestamp 1666464484
transform 1 0 40480 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_435
timestamp 1666464484
transform 1 0 41124 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_439
timestamp 1666464484
transform 1 0 41492 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_98_445
timestamp 1666464484
transform 1 0 42044 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_449
timestamp 1666464484
transform 1 0 42412 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_98_456
timestamp 1666464484
transform 1 0 43056 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_463
timestamp 1666464484
transform 1 0 43700 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_471
timestamp 1666464484
transform 1 0 44436 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1666464484
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_477
timestamp 1666464484
transform 1 0 44988 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_98_486
timestamp 1666464484
transform 1 0 45816 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_98_492
timestamp 1666464484
transform 1 0 46368 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_98_498
timestamp 1666464484
transform 1 0 46920 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_506
timestamp 1666464484
transform 1 0 47656 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_514
timestamp 1666464484
transform 1 0 48392 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_522
timestamp 1666464484
transform 1 0 49128 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_530
timestamp 1666464484
transform 1 0 49864 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_98_533
timestamp 1666464484
transform 1 0 50140 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_541
timestamp 1666464484
transform 1 0 50876 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_549
timestamp 1666464484
transform 1 0 51612 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_557
timestamp 1666464484
transform 1 0 52348 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_565
timestamp 1666464484
transform 1 0 53084 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_573
timestamp 1666464484
transform 1 0 53820 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_98_581
timestamp 1666464484
transform 1 0 54556 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_98_585
timestamp 1666464484
transform 1 0 54924 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1666464484
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_98_589
timestamp 1666464484
transform 1 0 55292 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_597
timestamp 1666464484
transform 1 0 56028 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_605
timestamp 1666464484
transform 1 0 56764 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_98_613
timestamp 1666464484
transform 1 0 57500 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_98_621
timestamp 1666464484
transform 1 0 58236 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_99_3
timestamp 1666464484
transform 1 0 1380 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_11
timestamp 1666464484
transform 1 0 2116 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_19
timestamp 1666464484
transform 1 0 2852 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_27
timestamp 1666464484
transform 1 0 3588 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_35
timestamp 1666464484
transform 1 0 4324 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_43
timestamp 1666464484
transform 1 0 5060 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_99_51
timestamp 1666464484
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1666464484
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_99_57
timestamp 1666464484
transform 1 0 6348 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_65
timestamp 1666464484
transform 1 0 7084 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_73
timestamp 1666464484
transform 1 0 7820 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_81
timestamp 1666464484
transform 1 0 8556 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_89
timestamp 1666464484
transform 1 0 9292 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_97
timestamp 1666464484
transform 1 0 10028 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_99_105
timestamp 1666464484
transform 1 0 10764 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_109
timestamp 1666464484
transform 1 0 11132 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1666464484
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_99_113
timestamp 1666464484
transform 1 0 11500 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_121
timestamp 1666464484
transform 1 0 12236 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_129
timestamp 1666464484
transform 1 0 12972 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_137
timestamp 1666464484
transform 1 0 13708 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_145
timestamp 1666464484
transform 1 0 14444 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_153
timestamp 1666464484
transform 1 0 15180 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_99_161
timestamp 1666464484
transform 1 0 15916 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_165
timestamp 1666464484
transform 1 0 16284 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1666464484
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_99_169
timestamp 1666464484
transform 1 0 16652 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_177
timestamp 1666464484
transform 1 0 17388 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_185
timestamp 1666464484
transform 1 0 18124 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_193
timestamp 1666464484
transform 1 0 18860 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_201
timestamp 1666464484
transform 1 0 19596 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_209
timestamp 1666464484
transform 1 0 20332 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_99_217
timestamp 1666464484
transform 1 0 21068 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_221
timestamp 1666464484
transform 1 0 21436 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1666464484
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_99_225
timestamp 1666464484
transform 1 0 21804 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_233
timestamp 1666464484
transform 1 0 22540 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_99_237
timestamp 1666464484
transform 1 0 22908 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_241
timestamp 1666464484
transform 1 0 23276 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_99_245
timestamp 1666464484
transform 1 0 23644 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_255
timestamp 1666464484
transform 1 0 24564 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_259
timestamp 1666464484
transform 1 0 24932 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_261
timestamp 1666464484
transform 1 0 25116 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_99_267
timestamp 1666464484
transform 1 0 25668 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_271
timestamp 1666464484
transform 1 0 26036 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_278
timestamp 1666464484
transform 1 0 26680 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_281
timestamp 1666464484
transform 1 0 26956 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_99_291
timestamp 1666464484
transform 1 0 27876 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_300
timestamp 1666464484
transform 1 0 28704 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_308
timestamp 1666464484
transform 1 0 29440 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_312
timestamp 1666464484
transform 1 0 29808 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_99_317
timestamp 1666464484
transform 1 0 30268 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_321
timestamp 1666464484
transform 1 0 30636 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_99_330
timestamp 1666464484
transform 1 0 31464 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_334
timestamp 1666464484
transform 1 0 31832 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_99_337
timestamp 1666464484
transform 1 0 32108 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_344
timestamp 1666464484
transform 1 0 32752 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_355
timestamp 1666464484
transform 1 0 33764 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_99_365
timestamp 1666464484
transform 1 0 34684 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_99_378
timestamp 1666464484
transform 1 0 35880 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_382
timestamp 1666464484
transform 1 0 36248 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_390
timestamp 1666464484
transform 1 0 36984 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_99_393
timestamp 1666464484
transform 1 0 37260 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_397
timestamp 1666464484
transform 1 0 37628 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_99_404
timestamp 1666464484
transform 1 0 38272 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_413
timestamp 1666464484
transform 1 0 39100 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_419
timestamp 1666464484
transform 1 0 39652 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_431
timestamp 1666464484
transform 1 0 40756 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_435
timestamp 1666464484
transform 1 0 41124 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_437
timestamp 1666464484
transform 1 0 41308 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_99_444
timestamp 1666464484
transform 1 0 41952 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_449
timestamp 1666464484
transform 1 0 42412 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_99_458
timestamp 1666464484
transform 1 0 43240 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_468
timestamp 1666464484
transform 1 0 44160 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_479
timestamp 1666464484
transform 1 0 45172 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_488
timestamp 1666464484
transform 1 0 46000 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_495
timestamp 1666464484
transform 1 0 46644 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_502
timestamp 1666464484
transform 1 0 47288 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_99_505
timestamp 1666464484
transform 1 0 47564 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_512
timestamp 1666464484
transform 1 0 48208 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_516
timestamp 1666464484
transform 1 0 48576 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_518
timestamp 1666464484
transform 1 0 48760 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_99_522
timestamp 1666464484
transform 1 0 49128 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_99_529
timestamp 1666464484
transform 1 0 49772 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_99_535
timestamp 1666464484
transform 1 0 50324 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_99_543
timestamp 1666464484
transform 1 0 51060 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_99_549
timestamp 1666464484
transform 1 0 51612 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_557
timestamp 1666464484
transform 1 0 52348 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1666464484
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_561
timestamp 1666464484
transform 1 0 52716 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_99_565
timestamp 1666464484
transform 1 0 53084 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_573
timestamp 1666464484
transform 1 0 53820 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_581
timestamp 1666464484
transform 1 0 54556 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_589
timestamp 1666464484
transform 1 0 55292 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_597
timestamp 1666464484
transform 1 0 56028 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_99_605
timestamp 1666464484
transform 1 0 56764 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_613
timestamp 1666464484
transform 1 0 57500 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1666464484
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_99_617
timestamp 1666464484
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_3
timestamp 1666464484
transform 1 0 1380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_11
timestamp 1666464484
transform 1 0 2116 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_19
timestamp 1666464484
transform 1 0 2852 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1666464484
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_100_29
timestamp 1666464484
transform 1 0 3772 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_37
timestamp 1666464484
transform 1 0 4508 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_100_42
timestamp 1666464484
transform 1 0 4968 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_50
timestamp 1666464484
transform 1 0 5704 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_55
timestamp 1666464484
transform 1 0 6164 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_100_62
timestamp 1666464484
transform 1 0 6808 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_70
timestamp 1666464484
transform 1 0 7544 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_100_78
timestamp 1666464484
transform 1 0 8280 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_82
timestamp 1666464484
transform 1 0 8648 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_100_85
timestamp 1666464484
transform 1 0 8924 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_93
timestamp 1666464484
transform 1 0 9660 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_100_101
timestamp 1666464484
transform 1 0 10396 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_105
timestamp 1666464484
transform 1 0 10764 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_107
timestamp 1666464484
transform 1 0 10948 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_100_110
timestamp 1666464484
transform 1 0 11224 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_100_117
timestamp 1666464484
transform 1 0 11868 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_125
timestamp 1666464484
transform 1 0 12604 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_100_133
timestamp 1666464484
transform 1 0 13340 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_137
timestamp 1666464484
transform 1 0 13708 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1666464484
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_141
timestamp 1666464484
transform 1 0 14076 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_143
timestamp 1666464484
transform 1 0 14260 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_100_147
timestamp 1666464484
transform 1 0 14628 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_155
timestamp 1666464484
transform 1 0 15364 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_163
timestamp 1666464484
transform 1 0 16100 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_171
timestamp 1666464484
transform 1 0 16836 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_173
timestamp 1666464484
transform 1 0 17020 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_100_177
timestamp 1666464484
transform 1 0 17388 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_185
timestamp 1666464484
transform 1 0 18124 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_193
timestamp 1666464484
transform 1 0 18860 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1666464484
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_100_197
timestamp 1666464484
transform 1 0 19228 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_201
timestamp 1666464484
transform 1 0 19596 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_203
timestamp 1666464484
transform 1 0 19780 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_100_207
timestamp 1666464484
transform 1 0 20148 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_215
timestamp 1666464484
transform 1 0 20884 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_220
timestamp 1666464484
transform 1 0 21344 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_228
timestamp 1666464484
transform 1 0 22080 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_232
timestamp 1666464484
transform 1 0 22448 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_234
timestamp 1666464484
transform 1 0 22632 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_100_238
timestamp 1666464484
transform 1 0 23000 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_250
timestamp 1666464484
transform 1 0 24104 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_253
timestamp 1666464484
transform 1 0 24380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_257
timestamp 1666464484
transform 1 0 24748 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_259
timestamp 1666464484
transform 1 0 24932 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_100_268
timestamp 1666464484
transform 1 0 25760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_276
timestamp 1666464484
transform 1 0 26496 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_100_280
timestamp 1666464484
transform 1 0 26864 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_291
timestamp 1666464484
transform 1 0 27876 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_295
timestamp 1666464484
transform 1 0 28244 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_297
timestamp 1666464484
transform 1 0 28428 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_306
timestamp 1666464484
transform 1 0 29256 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_309
timestamp 1666464484
transform 1 0 29532 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_320
timestamp 1666464484
transform 1 0 30544 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_324
timestamp 1666464484
transform 1 0 30912 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_329
timestamp 1666464484
transform 1 0 31372 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_341
timestamp 1666464484
transform 1 0 32476 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_351
timestamp 1666464484
transform 1 0 33396 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_361
timestamp 1666464484
transform 1 0 34316 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1666464484
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_100_365
timestamp 1666464484
transform 1 0 34684 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_377
timestamp 1666464484
transform 1 0 35788 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_381
timestamp 1666464484
transform 1 0 36156 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_100_392
timestamp 1666464484
transform 1 0 37168 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_400
timestamp 1666464484
transform 1 0 37904 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_100_408
timestamp 1666464484
transform 1 0 38640 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_416
timestamp 1666464484
transform 1 0 39376 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_421
timestamp 1666464484
transform 1 0 39836 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_430
timestamp 1666464484
transform 1 0 40664 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_442
timestamp 1666464484
transform 1 0 41768 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_449
timestamp 1666464484
transform 1 0 42412 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_455
timestamp 1666464484
transform 1 0 42964 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_469
timestamp 1666464484
transform 1 0 44252 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_473
timestamp 1666464484
transform 1 0 44620 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1666464484
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_477
timestamp 1666464484
transform 1 0 44988 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_482
timestamp 1666464484
transform 1 0 45448 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_489
timestamp 1666464484
transform 1 0 46092 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_496
timestamp 1666464484
transform 1 0 46736 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_503
timestamp 1666464484
transform 1 0 47380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_510
timestamp 1666464484
transform 1 0 48024 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_524
timestamp 1666464484
transform 1 0 49312 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_530
timestamp 1666464484
transform 1 0 49864 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_533
timestamp 1666464484
transform 1 0 50140 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_538
timestamp 1666464484
transform 1 0 50600 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_545
timestamp 1666464484
transform 1 0 51244 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_552
timestamp 1666464484
transform 1 0 51888 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_559
timestamp 1666464484
transform 1 0 52532 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_563
timestamp 1666464484
transform 1 0 52900 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_100_567
timestamp 1666464484
transform 1 0 53268 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_100_574
timestamp 1666464484
transform 1 0 53912 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_100_580
timestamp 1666464484
transform 1 0 54464 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_589
timestamp 1666464484
transform 1 0 55292 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_100_594
timestamp 1666464484
transform 1 0 55752 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_100_600
timestamp 1666464484
transform 1 0 56304 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_608
timestamp 1666464484
transform 1 0 57040 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_100_616
timestamp 1666464484
transform 1 0 57776 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_624
timestamp 1666464484
transform 1 0 58512 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_101_3
timestamp 1666464484
transform 1 0 1380 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_101_11
timestamp 1666464484
transform 1 0 2116 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_101_19
timestamp 1666464484
transform 1 0 2852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_23
timestamp 1666464484
transform 1 0 3220 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_26
timestamp 1666464484
transform 1 0 3496 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_29
timestamp 1666464484
transform 1 0 3772 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_101_35
timestamp 1666464484
transform 1 0 4324 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_43
timestamp 1666464484
transform 1 0 5060 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_48
timestamp 1666464484
transform 1 0 5520 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1666464484
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_101_57
timestamp 1666464484
transform 1 0 6348 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_101_68
timestamp 1666464484
transform 1 0 7360 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_75
timestamp 1666464484
transform 1 0 8004 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_82
timestamp 1666464484
transform 1 0 8648 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_85
timestamp 1666464484
transform 1 0 8924 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_92
timestamp 1666464484
transform 1 0 9568 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_96
timestamp 1666464484
transform 1 0 9936 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_100
timestamp 1666464484
transform 1 0 10304 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_108
timestamp 1666464484
transform 1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_113
timestamp 1666464484
transform 1 0 11500 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_117
timestamp 1666464484
transform 1 0 11868 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_123
timestamp 1666464484
transform 1 0 12420 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_130
timestamp 1666464484
transform 1 0 13064 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_138
timestamp 1666464484
transform 1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_101_141
timestamp 1666464484
transform 1 0 14076 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_101_153
timestamp 1666464484
transform 1 0 15180 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_157
timestamp 1666464484
transform 1 0 15548 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_162
timestamp 1666464484
transform 1 0 16008 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_166
timestamp 1666464484
transform 1 0 16376 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_169
timestamp 1666464484
transform 1 0 16652 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_175
timestamp 1666464484
transform 1 0 17204 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_183
timestamp 1666464484
transform 1 0 17940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_187
timestamp 1666464484
transform 1 0 18308 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_192
timestamp 1666464484
transform 1 0 18768 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_197
timestamp 1666464484
transform 1 0 19228 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_203
timestamp 1666464484
transform 1 0 19780 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_207
timestamp 1666464484
transform 1 0 20148 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_213
timestamp 1666464484
transform 1 0 20700 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_217
timestamp 1666464484
transform 1 0 21068 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_222
timestamp 1666464484
transform 1 0 21528 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_225
timestamp 1666464484
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_233
timestamp 1666464484
transform 1 0 22540 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_241
timestamp 1666464484
transform 1 0 23276 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_250
timestamp 1666464484
transform 1 0 24104 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_253
timestamp 1666464484
transform 1 0 24380 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_101_260
timestamp 1666464484
transform 1 0 25024 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_268
timestamp 1666464484
transform 1 0 25760 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_273
timestamp 1666464484
transform 1 0 26220 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_277
timestamp 1666464484
transform 1 0 26588 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1666464484
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_281
timestamp 1666464484
transform 1 0 26956 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_283
timestamp 1666464484
transform 1 0 27140 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_288
timestamp 1666464484
transform 1 0 27600 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_295
timestamp 1666464484
transform 1 0 28244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_303
timestamp 1666464484
transform 1 0 28980 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_307
timestamp 1666464484
transform 1 0 29348 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_309
timestamp 1666464484
transform 1 0 29532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_313
timestamp 1666464484
transform 1 0 29900 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_315
timestamp 1666464484
transform 1 0 30084 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_319
timestamp 1666464484
transform 1 0 30452 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_326
timestamp 1666464484
transform 1 0 31096 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_334
timestamp 1666464484
transform 1 0 31832 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_337
timestamp 1666464484
transform 1 0 32108 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_349
timestamp 1666464484
transform 1 0 33212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_359
timestamp 1666464484
transform 1 0 34132 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_363
timestamp 1666464484
transform 1 0 34500 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_365
timestamp 1666464484
transform 1 0 34684 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_369
timestamp 1666464484
transform 1 0 35052 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_375
timestamp 1666464484
transform 1 0 35604 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_389
timestamp 1666464484
transform 1 0 36892 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1666464484
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_393
timestamp 1666464484
transform 1 0 37260 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_405
timestamp 1666464484
transform 1 0 38364 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_412
timestamp 1666464484
transform 1 0 39008 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_418
timestamp 1666464484
transform 1 0 39560 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_421
timestamp 1666464484
transform 1 0 39836 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_433
timestamp 1666464484
transform 1 0 40940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_443
timestamp 1666464484
transform 1 0 41860 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1666464484
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_449
timestamp 1666464484
transform 1 0 42412 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_453
timestamp 1666464484
transform 1 0 42780 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_464
timestamp 1666464484
transform 1 0 43792 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_474
timestamp 1666464484
transform 1 0 44712 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_477
timestamp 1666464484
transform 1 0 44988 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_481
timestamp 1666464484
transform 1 0 45356 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_483
timestamp 1666464484
transform 1 0 45540 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_488
timestamp 1666464484
transform 1 0 46000 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_495
timestamp 1666464484
transform 1 0 46644 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_502
timestamp 1666464484
transform 1 0 47288 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_505
timestamp 1666464484
transform 1 0 47564 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_517
timestamp 1666464484
transform 1 0 48668 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_524
timestamp 1666464484
transform 1 0 49312 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_530
timestamp 1666464484
transform 1 0 49864 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1666464484
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_545
timestamp 1666464484
transform 1 0 51244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_553
timestamp 1666464484
transform 1 0 51980 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_557
timestamp 1666464484
transform 1 0 52348 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1666464484
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_561
timestamp 1666464484
transform 1 0 52716 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_569
timestamp 1666464484
transform 1 0 53452 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_573
timestamp 1666464484
transform 1 0 53820 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_101_578
timestamp 1666464484
transform 1 0 54280 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_585
timestamp 1666464484
transform 1 0 54924 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_587
timestamp 1666464484
transform 1 0 55108 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_589
timestamp 1666464484
transform 1 0 55292 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_101_595
timestamp 1666464484
transform 1 0 55844 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_602
timestamp 1666464484
transform 1 0 56488 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_101_609
timestamp 1666464484
transform 1 0 57132 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_101_613
timestamp 1666464484
transform 1 0 57500 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1666464484
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_101_617
timestamp 1666464484
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1666464484
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1666464484
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1666464484
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1666464484
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1666464484
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1666464484
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1666464484
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1666464484
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1666464484
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1666464484
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1666464484
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1666464484
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1666464484
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1666464484
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1666464484
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1666464484
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1666464484
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1666464484
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1666464484
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1666464484
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1666464484
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1666464484
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1666464484
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1666464484
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1666464484
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1666464484
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1666464484
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1666464484
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1666464484
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1666464484
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1666464484
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1666464484
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1666464484
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1666464484
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1666464484
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1666464484
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1666464484
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1666464484
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1666464484
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1666464484
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1666464484
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1666464484
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1666464484
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1666464484
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1666464484
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1666464484
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1666464484
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1666464484
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1666464484
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1666464484
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1666464484
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1666464484
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1666464484
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1666464484
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1666464484
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1666464484
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1666464484
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1666464484
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1666464484
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1666464484
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1666464484
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1666464484
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1666464484
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1666464484
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1666464484
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1666464484
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1666464484
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1666464484
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1666464484
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1666464484
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1666464484
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1666464484
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1666464484
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1666464484
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1666464484
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1666464484
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1666464484
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1666464484
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1666464484
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1666464484
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1666464484
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1666464484
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1666464484
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1666464484
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1666464484
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1666464484
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1666464484
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1666464484
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1666464484
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1666464484
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1666464484
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1666464484
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1666464484
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1666464484
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1666464484
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1666464484
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1666464484
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1666464484
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1666464484
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1666464484
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1666464484
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1666464484
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1666464484
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1666464484
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1666464484
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1666464484
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1666464484
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1666464484
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1666464484
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1666464484
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1666464484
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1666464484
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1666464484
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1666464484
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1666464484
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1666464484
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1666464484
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1666464484
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1666464484
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1666464484
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1666464484
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1666464484
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1666464484
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1666464484
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1666464484
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1666464484
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1666464484
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1666464484
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1666464484
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1666464484
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1666464484
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1666464484
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1666464484
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1666464484
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1666464484
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1666464484
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1666464484
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1666464484
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1666464484
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1666464484
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1666464484
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1666464484
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1666464484
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1666464484
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1666464484
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1666464484
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1666464484
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1666464484
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1666464484
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1666464484
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1666464484
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1666464484
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1666464484
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1666464484
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1666464484
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1666464484
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1666464484
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1666464484
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1666464484
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1666464484
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1666464484
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1666464484
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1666464484
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1666464484
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1666464484
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1666464484
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1666464484
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1666464484
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1666464484
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1666464484
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1666464484
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1666464484
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1666464484
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1666464484
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1666464484
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1666464484
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1666464484
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1666464484
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1666464484
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1666464484
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1666464484
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1666464484
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1666464484
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1666464484
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1666464484
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1666464484
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1666464484
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1666464484
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1666464484
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1666464484
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1666464484
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1666464484
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1666464484
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1666464484
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1666464484
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1666464484
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1666464484
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1666464484
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1666464484
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1666464484
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1666464484
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1666464484
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1666464484
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1666464484
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1666464484
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1666464484
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1666464484
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1666464484
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1666464484
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1666464484
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1666464484
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1666464484
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1666464484
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1666464484
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1666464484
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1666464484
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1666464484
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1666464484
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1666464484
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1666464484
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1666464484
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1666464484
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1666464484
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1666464484
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1666464484
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1666464484
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1666464484
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1666464484
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1666464484
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1666464484
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1666464484
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1666464484
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1666464484
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1666464484
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1666464484
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1666464484
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1666464484
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1666464484
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1666464484
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1666464484
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1666464484
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1666464484
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1666464484
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1666464484
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1666464484
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1666464484
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1666464484
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1666464484
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1666464484
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1666464484
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1666464484
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1666464484
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1666464484
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1666464484
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1666464484
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1666464484
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1666464484
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1666464484
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1666464484
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1666464484
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1666464484
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1666464484
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1666464484
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1666464484
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1666464484
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1666464484
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1666464484
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1666464484
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1666464484
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1666464484
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1666464484
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1666464484
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1666464484
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1666464484
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1666464484
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1666464484
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1666464484
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1666464484
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1666464484
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1666464484
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1666464484
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1666464484
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1666464484
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1666464484
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1666464484
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1666464484
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1666464484
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1666464484
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1666464484
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1666464484
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1666464484
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1666464484
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1666464484
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1666464484
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1666464484
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1666464484
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1666464484
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1666464484
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1666464484
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1666464484
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1666464484
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1666464484
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1666464484
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1666464484
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1666464484
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1666464484
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1666464484
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1666464484
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1666464484
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1666464484
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1666464484
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1666464484
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1666464484
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1666464484
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1666464484
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1666464484
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1666464484
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1666464484
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1666464484
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1666464484
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1666464484
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1666464484
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1666464484
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1666464484
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1666464484
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1666464484
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1666464484
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1666464484
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1666464484
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1666464484
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1666464484
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1666464484
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1666464484
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1666464484
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1666464484
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1666464484
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1666464484
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1666464484
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1666464484
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1666464484
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1666464484
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1666464484
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1666464484
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1666464484
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1666464484
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1666464484
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1666464484
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1666464484
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1666464484
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1666464484
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1666464484
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1666464484
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1666464484
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1666464484
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1666464484
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1666464484
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1666464484
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1666464484
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1666464484
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1666464484
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1666464484
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1666464484
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1666464484
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1666464484
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1666464484
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1666464484
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1666464484
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1666464484
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1666464484
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1666464484
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1666464484
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1666464484
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1666464484
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1666464484
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1666464484
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1666464484
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1666464484
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1666464484
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1666464484
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1666464484
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1666464484
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1666464484
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1666464484
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1666464484
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1666464484
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1666464484
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1666464484
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1666464484
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1666464484
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1666464484
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1666464484
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1666464484
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1666464484
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1666464484
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1666464484
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1666464484
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1666464484
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1666464484
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1666464484
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1666464484
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1666464484
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1666464484
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1666464484
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1666464484
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1666464484
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1666464484
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1666464484
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1666464484
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1666464484
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1666464484
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1666464484
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1666464484
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1666464484
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1666464484
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1666464484
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1666464484
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1666464484
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1666464484
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1666464484
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1666464484
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1666464484
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1666464484
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1666464484
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1666464484
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1666464484
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1666464484
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1666464484
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1666464484
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1666464484
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1666464484
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1666464484
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1666464484
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1666464484
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1666464484
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1666464484
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1666464484
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1666464484
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1666464484
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1666464484
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1666464484
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1666464484
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1666464484
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1666464484
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1666464484
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1666464484
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1666464484
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1666464484
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1666464484
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1666464484
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1666464484
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1666464484
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1666464484
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1666464484
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1666464484
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1666464484
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1666464484
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1666464484
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1666464484
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1666464484
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1666464484
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1666464484
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1666464484
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1666464484
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1666464484
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1666464484
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1666464484
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1666464484
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1666464484
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1666464484
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1666464484
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1666464484
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1666464484
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1666464484
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1666464484
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1666464484
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1666464484
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1666464484
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1666464484
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1666464484
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1666464484
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1666464484
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1666464484
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1666464484
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1666464484
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1666464484
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1666464484
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1666464484
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1666464484
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1666464484
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1666464484
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1666464484
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1666464484
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1666464484
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1666464484
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1666464484
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1666464484
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1666464484
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1666464484
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1666464484
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1666464484
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1666464484
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1666464484
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1666464484
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1666464484
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1666464484
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1666464484
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1666464484
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1666464484
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1666464484
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1666464484
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1666464484
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1666464484
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1666464484
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1666464484
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1666464484
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1666464484
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1666464484
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1666464484
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1666464484
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1666464484
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1666464484
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1666464484
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1666464484
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1666464484
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1666464484
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1666464484
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1666464484
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1666464484
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1666464484
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1666464484
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1666464484
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1666464484
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1666464484
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1666464484
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1666464484
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1666464484
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1666464484
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1666464484
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1666464484
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1666464484
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1666464484
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1666464484
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1666464484
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1666464484
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1666464484
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1666464484
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1666464484
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1666464484
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1666464484
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1666464484
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1666464484
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1666464484
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1666464484
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1666464484
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1666464484
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1666464484
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1666464484
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1666464484
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1666464484
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1666464484
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1666464484
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1666464484
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1666464484
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1666464484
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1666464484
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1666464484
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1666464484
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1666464484
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1666464484
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1666464484
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1666464484
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1666464484
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1666464484
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1666464484
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1666464484
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1666464484
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1666464484
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1666464484
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1666464484
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1666464484
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1666464484
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1666464484
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1666464484
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1666464484
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1666464484
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1666464484
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1666464484
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1666464484
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1666464484
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1666464484
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1666464484
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1666464484
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1666464484
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1666464484
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1666464484
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1666464484
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1666464484
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1666464484
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1666464484
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1666464484
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1666464484
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1666464484
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1666464484
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1666464484
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1666464484
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1666464484
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1666464484
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1666464484
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1666464484
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1666464484
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1666464484
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1666464484
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1666464484
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1666464484
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1666464484
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1666464484
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1666464484
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1666464484
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1666464484
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1666464484
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1666464484
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1666464484
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1666464484
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1666464484
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1666464484
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1666464484
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1666464484
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1666464484
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1666464484
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1666464484
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1666464484
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1666464484
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1666464484
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1666464484
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1666464484
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1666464484
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1666464484
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1666464484
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1666464484
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1666464484
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1666464484
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1666464484
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1666464484
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1666464484
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1666464484
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1666464484
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1666464484
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1666464484
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1666464484
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1666464484
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1666464484
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1666464484
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1666464484
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1666464484
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1666464484
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1666464484
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1666464484
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1666464484
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1666464484
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1666464484
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1666464484
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1666464484
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1666464484
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1666464484
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1666464484
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1666464484
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1666464484
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1666464484
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1666464484
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1666464484
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1666464484
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1666464484
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1666464484
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1666464484
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1666464484
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1666464484
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1666464484
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1666464484
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1666464484
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1666464484
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1666464484
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1666464484
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1666464484
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1666464484
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1666464484
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1666464484
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1666464484
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1666464484
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1666464484
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1666464484
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1666464484
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1666464484
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1666464484
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1666464484
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1666464484
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1666464484
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1666464484
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1666464484
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1666464484
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1666464484
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1666464484
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1666464484
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1666464484
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1666464484
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1666464484
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1666464484
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1666464484
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1666464484
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1666464484
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1666464484
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1666464484
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1666464484
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1666464484
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1666464484
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1666464484
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1666464484
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1666464484
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1666464484
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1666464484
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1666464484
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1666464484
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1666464484
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1666464484
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1666464484
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1666464484
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1666464484
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1666464484
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1666464484
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1666464484
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1666464484
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1666464484
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1666464484
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1666464484
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1666464484
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1666464484
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1666464484
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1666464484
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1666464484
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1666464484
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1666464484
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1666464484
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1666464484
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1666464484
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1666464484
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1666464484
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1666464484
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1666464484
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1666464484
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1666464484
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1666464484
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1666464484
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1666464484
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1666464484
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1666464484
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1666464484
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1666464484
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1666464484
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1666464484
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1666464484
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1666464484
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1666464484
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1666464484
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1666464484
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1666464484
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1666464484
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1666464484
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1666464484
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1666464484
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1666464484
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1666464484
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1666464484
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1666464484
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1666464484
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1666464484
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1666464484
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1666464484
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1666464484
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1666464484
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1666464484
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1666464484
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1666464484
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1666464484
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1666464484
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1666464484
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1666464484
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1666464484
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1666464484
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1666464484
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1666464484
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1666464484
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1666464484
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1666464484
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1666464484
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1666464484
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1666464484
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1666464484
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1666464484
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1666464484
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1666464484
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1666464484
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1666464484
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1666464484
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1666464484
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1666464484
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1666464484
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1666464484
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1666464484
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1666464484
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1666464484
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1666464484
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1666464484
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1666464484
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1666464484
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1666464484
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1666464484
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1666464484
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1666464484
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1666464484
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1666464484
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1666464484
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1666464484
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1666464484
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1666464484
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1666464484
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1666464484
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1666464484
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1666464484
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1666464484
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1666464484
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1666464484
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1666464484
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1666464484
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1666464484
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1666464484
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1666464484
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1666464484
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1666464484
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1666464484
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1666464484
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1666464484
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1666464484
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1666464484
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1666464484
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1666464484
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1666464484
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1666464484
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1666464484
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1666464484
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1666464484
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1666464484
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1666464484
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1666464484
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1666464484
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1666464484
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1666464484
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1666464484
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1666464484
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1666464484
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1666464484
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1666464484
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1666464484
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1666464484
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1666464484
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1666464484
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1666464484
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1666464484
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1666464484
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1666464484
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1666464484
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1666464484
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1666464484
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1666464484
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1666464484
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1666464484
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1666464484
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1666464484
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1666464484
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1666464484
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1666464484
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1666464484
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1666464484
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1666464484
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1666464484
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1666464484
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1666464484
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1666464484
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1666464484
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1666464484
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1666464484
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1666464484
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1666464484
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1666464484
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1666464484
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1666464484
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1666464484
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1666464484
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1666464484
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1666464484
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1666464484
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1666464484
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1666464484
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1666464484
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1666464484
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1666464484
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1666464484
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1666464484
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1666464484
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1666464484
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1666464484
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1666464484
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1666464484
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1666464484
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1666464484
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1666464484
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1666464484
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1666464484
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1666464484
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1666464484
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1666464484
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1666464484
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1666464484
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1666464484
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1666464484
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1666464484
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1666464484
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1666464484
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1666464484
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1666464484
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1666464484
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1666464484
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1666464484
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1666464484
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1666464484
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1666464484
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1666464484
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1666464484
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1666464484
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1666464484
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1666464484
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1666464484
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1666464484
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1666464484
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1666464484
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1666464484
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1666464484
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1666464484
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1666464484
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1666464484
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1666464484
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1666464484
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1666464484
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1666464484
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1666464484
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1666464484
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1666464484
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1666464484
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1666464484
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1666464484
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1666464484
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1666464484
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1666464484
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1666464484
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1666464484
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1666464484
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1666464484
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1666464484
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1666464484
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1666464484
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1666464484
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1666464484
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1666464484
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1666464484
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1666464484
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1666464484
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1666464484
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1666464484
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1666464484
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1666464484
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1666464484
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1666464484
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1666464484
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1666464484
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1666464484
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1666464484
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1666464484
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1666464484
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1666464484
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1666464484
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1666464484
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1666464484
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1666464484
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1666464484
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1666464484
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1666464484
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1666464484
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1666464484
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1666464484
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1666464484
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1666464484
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1666464484
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1666464484
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1666464484
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1666464484
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1666464484
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1666464484
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1666464484
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1666464484
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1666464484
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1666464484
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1666464484
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1666464484
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1666464484
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1666464484
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1666464484
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1666464484
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1666464484
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1666464484
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1666464484
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1666464484
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1666464484
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1666464484
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1666464484
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1666464484
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1666464484
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1666464484
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1666464484
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1666464484
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1666464484
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1666464484
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1666464484
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1666464484
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1666464484
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1666464484
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1666464484
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1666464484
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1666464484
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1666464484
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1666464484
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1666464484
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1666464484
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1666464484
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1666464484
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1666464484
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1666464484
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1666464484
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1666464484
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1666464484
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1666464484
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1666464484
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1666464484
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1666464484
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1666464484
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1666464484
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1666464484
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1666464484
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1666464484
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1666464484
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1666464484
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1666464484
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1666464484
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1666464484
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1666464484
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1666464484
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1666464484
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1666464484
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1666464484
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1666464484
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1666464484
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1666464484
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1666464484
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1666464484
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1666464484
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1666464484
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1666464484
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1666464484
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1666464484
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1666464484
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1666464484
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1666464484
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1666464484
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1666464484
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1666464484
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1666464484
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1666464484
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1666464484
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1666464484
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1666464484
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1666464484
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1666464484
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1666464484
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1666464484
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1666464484
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1666464484
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1666464484
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1666464484
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1666464484
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1666464484
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1666464484
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1666464484
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1666464484
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1666464484
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1666464484
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1666464484
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1666464484
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1666464484
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1666464484
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1666464484
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1666464484
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1666464484
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1666464484
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1666464484
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1666464484
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1666464484
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1666464484
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1666464484
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1666464484
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1666464484
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1666464484
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1666464484
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1666464484
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1666464484
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1666464484
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1666464484
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1666464484
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1666464484
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1666464484
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1666464484
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1666464484
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1666464484
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1666464484
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1666464484
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1666464484
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1666464484
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1666464484
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1666464484
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1666464484
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1666464484
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1666464484
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1666464484
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1666464484
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1666464484
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1666464484
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1666464484
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1666464484
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1666464484
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1666464484
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1666464484
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1666464484
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1666464484
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1666464484
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1666464484
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1666464484
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1666464484
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1666464484
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1666464484
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1666464484
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1666464484
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1666464484
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1666464484
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1666464484
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1666464484
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1666464484
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1666464484
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1666464484
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1666464484
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1666464484
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1666464484
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1666464484
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1666464484
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1666464484
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1666464484
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1666464484
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1666464484
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1666464484
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1666464484
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1666464484
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1666464484
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1666464484
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1666464484
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1666464484
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1666464484
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1666464484
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1666464484
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1666464484
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1666464484
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1666464484
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1666464484
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1666464484
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1666464484
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1666464484
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1666464484
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1666464484
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1666464484
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1666464484
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1666464484
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1666464484
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1666464484
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1666464484
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1666464484
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1666464484
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1666464484
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1666464484
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1666464484
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1666464484
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1666464484
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1666464484
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1666464484
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1666464484
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1666464484
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1666464484
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1666464484
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1666464484
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1666464484
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1666464484
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1666464484
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1666464484
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1666464484
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1666464484
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1666464484
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1666464484
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1666464484
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1666464484
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1666464484
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1666464484
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1666464484
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1666464484
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1666464484
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1666464484
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1666464484
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1666464484
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1666464484
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1666464484
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1666464484
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1666464484
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1666464484
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1666464484
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1666464484
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1666464484
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1666464484
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1666464484
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1666464484
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1666464484
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1666464484
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1666464484
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1666464484
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1666464484
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1666464484
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1666464484
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1666464484
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1666464484
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1666464484
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1666464484
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1666464484
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1666464484
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1666464484
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1666464484
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1666464484
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1666464484
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1666464484
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1666464484
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1666464484
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1666464484
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1666464484
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1666464484
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1666464484
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1666464484
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1666464484
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1666464484
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1666464484
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1666464484
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1666464484
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1666464484
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1666464484
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1666464484
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1666464484
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1666464484
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1666464484
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1666464484
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1666464484
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1666464484
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1666464484
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1666464484
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1666464484
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1666464484
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1666464484
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1666464484
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1666464484
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1666464484
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1666464484
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1666464484
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1666464484
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1666464484
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1666464484
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1666464484
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1666464484
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1666464484
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1666464484
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1666464484
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1666464484
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1666464484
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1666464484
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1666464484
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1666464484
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1666464484
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1666464484
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1666464484
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1666464484
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1666464484
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1666464484
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1666464484
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1666464484
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1666464484
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1666464484
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1666464484
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1666464484
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1666464484
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1666464484
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1666464484
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1666464484
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1666464484
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1666464484
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1666464484
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1666464484
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1666464484
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1666464484
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1666464484
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1666464484
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1666464484
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1666464484
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1666464484
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1666464484
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1666464484
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1666464484
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1666464484
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1666464484
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1666464484
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1666464484
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1666464484
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1666464484
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1666464484
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1666464484
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1666464484
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1666464484
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1666464484
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1666464484
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1666464484
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _157_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 26956 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 24012 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _159_
timestamp 1666464484
transform 1 0 32752 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1666464484
transform 1 0 38088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1666464484
transform -1 0 36432 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1666464484
transform -1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _163_
timestamp 1666464484
transform -1 0 37444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1666464484
transform -1 0 37720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1666464484
transform -1 0 35880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1666464484
transform -1 0 35144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _167_
timestamp 1666464484
transform 1 0 33672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1666464484
transform -1 0 35144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_
timestamp 1666464484
transform -1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _170_
timestamp 1666464484
transform 1 0 29716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _171_
timestamp 1666464484
transform -1 0 31372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _172_
timestamp 1666464484
transform 1 0 30452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1666464484
transform 1 0 25760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174_
timestamp 1666464484
transform 1 0 34960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1666464484
transform -1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _176_
timestamp 1666464484
transform -1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1666464484
transform -1 0 29992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp 1666464484
transform 1 0 28980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1666464484
transform 1 0 24104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1666464484
transform -1 0 24104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _181_
timestamp 1666464484
transform 1 0 27232 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1666464484
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp 1666464484
transform 1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1666464484
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1666464484
transform 1 0 27784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp 1666464484
transform 1 0 26404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1666464484
transform 1 0 26680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1666464484
transform 1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp 1666464484
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp 1666464484
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1666464484
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _192_
timestamp 1666464484
transform -1 0 25576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _193_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35880 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _194_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 35052 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _195_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35512 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _196_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30360 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _197_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 34868 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _198_
timestamp 1666464484
transform -1 0 35420 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _199_
timestamp 1666464484
transform -1 0 29808 0 -1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _200_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _201_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _202_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32844 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _203_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31740 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _204_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34040 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1666464484
transform 1 0 31924 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _206_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30268 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _207_
timestamp 1666464484
transform -1 0 30360 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _208_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30360 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _209_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 34408 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _210_
timestamp 1666464484
transform -1 0 28060 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _211_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 29072 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _212_
timestamp 1666464484
transform -1 0 28704 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _213_
timestamp 1666464484
transform -1 0 46000 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _214_
timestamp 1666464484
transform 1 0 45172 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _215_
timestamp 1666464484
transform -1 0 45172 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _216_
timestamp 1666464484
transform -1 0 39468 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _217_
timestamp 1666464484
transform -1 0 44252 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _218_
timestamp 1666464484
transform -1 0 44344 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _219_
timestamp 1666464484
transform -1 0 39652 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _220_
timestamp 1666464484
transform -1 0 43240 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _221_
timestamp 1666464484
transform -1 0 43332 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp 1666464484
transform -1 0 43148 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _223_
timestamp 1666464484
transform 1 0 40756 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1666464484
transform -1 0 42504 0 1 53312
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _225_
timestamp 1666464484
transform 1 0 41676 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _226_
timestamp 1666464484
transform -1 0 39100 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _227_
timestamp 1666464484
transform -1 0 38548 0 1 54400
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _228_
timestamp 1666464484
transform -1 0 38824 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _229_
timestamp 1666464484
transform -1 0 44436 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _230_
timestamp 1666464484
transform -1 0 39376 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _231_
timestamp 1666464484
transform 1 0 37996 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _232_
timestamp 1666464484
transform -1 0 35604 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_2  _233_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 35788 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _234_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 29072 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _235_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 27232 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1666464484
transform -1 0 32752 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _237_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 31740 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _238_
timestamp 1666464484
transform 1 0 32844 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _239_
timestamp 1666464484
transform 1 0 30820 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1666464484
transform -1 0 39284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _241_
timestamp 1666464484
transform 1 0 41032 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _242_
timestamp 1666464484
transform 1 0 41308 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _243_
timestamp 1666464484
transform 1 0 40020 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _244_
timestamp 1666464484
transform 1 0 23644 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _245_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 23828 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _246_
timestamp 1666464484
transform -1 0 25024 0 -1 57664
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1666464484
transform 1 0 23368 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _248_
timestamp 1666464484
transform -1 0 24104 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _249_
timestamp 1666464484
transform -1 0 33212 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _250_
timestamp 1666464484
transform 1 0 32292 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _251_
timestamp 1666464484
transform 1 0 34132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _252_
timestamp 1666464484
transform 1 0 33120 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _253_
timestamp 1666464484
transform 1 0 32936 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _254_
timestamp 1666464484
transform -1 0 41860 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 1666464484
transform 1 0 40940 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _256_
timestamp 1666464484
transform -1 0 43056 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _257_
timestamp 1666464484
transform 1 0 42596 0 -1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _258_
timestamp 1666464484
transform 1 0 41400 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _259_
timestamp 1666464484
transform -1 0 25760 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1666464484
transform 1 0 24656 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _261_
timestamp 1666464484
transform 1 0 25208 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1666464484
transform -1 0 25760 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _263_
timestamp 1666464484
transform -1 0 25760 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1666464484
transform 1 0 32016 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _265_
timestamp 1666464484
transform -1 0 32752 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _266_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 30176 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _267_
timestamp 1666464484
transform -1 0 31372 0 -1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _268_
timestamp 1666464484
transform 1 0 30820 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 31648 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _270_
timestamp 1666464484
transform -1 0 44160 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _271_
timestamp 1666464484
transform -1 0 42044 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _272_
timestamp 1666464484
transform 1 0 38916 0 1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _273_
timestamp 1666464484
transform -1 0 40480 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _274_
timestamp 1666464484
transform 1 0 40020 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _275_
timestamp 1666464484
transform -1 0 40756 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _276_
timestamp 1666464484
transform 1 0 26220 0 -1 56576
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _277_
timestamp 1666464484
transform 1 0 26404 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1666464484
transform 1 0 26680 0 1 55488
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _279_
timestamp 1666464484
transform -1 0 27416 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _280_
timestamp 1666464484
transform -1 0 27876 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _281_
timestamp 1666464484
transform 1 0 29072 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _282_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 28888 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _283_
timestamp 1666464484
transform -1 0 28888 0 -1 54400
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 26864 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _285_
timestamp 1666464484
transform 1 0 33764 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1666464484
transform 1 0 33580 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _287_
timestamp 1666464484
transform -1 0 28244 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _288_
timestamp 1666464484
transform 1 0 38088 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _289_
timestamp 1666464484
transform -1 0 38272 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _290_
timestamp 1666464484
transform 1 0 36524 0 1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _291_
timestamp 1666464484
transform 1 0 44160 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 43332 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _293_
timestamp 1666464484
transform 1 0 36432 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _294_
timestamp 1666464484
transform 1 0 36248 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 30544 0 1 56576
box -38 -48 866 592
use sky130_fd_sc_hd__o32a_1  _296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 28520 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _519__194 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform -1 0 25668 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 25024 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _520__195
timestamp 1666464484
transform 1 0 24472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _520_
timestamp 1666464484
transform 1 0 24748 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _521_
timestamp 1666464484
transform 1 0 25024 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _521__196
timestamp 1666464484
transform 1 0 22172 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _522__197
timestamp 1666464484
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _522_
timestamp 1666464484
transform 1 0 24748 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _523__198
timestamp 1666464484
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _523_
timestamp 1666464484
transform 1 0 26588 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _524__199
timestamp 1666464484
transform 1 0 26404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _524_
timestamp 1666464484
transform 1 0 27140 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _525__200
timestamp 1666464484
transform -1 0 28244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _525_
timestamp 1666464484
transform 1 0 27324 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _526__201
timestamp 1666464484
transform -1 0 27600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _526_
timestamp 1666464484
transform 1 0 27324 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _527__202
timestamp 1666464484
transform 1 0 25300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _527_
timestamp 1666464484
transform 1 0 27600 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _528__203
timestamp 1666464484
transform 1 0 24104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _528_
timestamp 1666464484
transform 1 0 27324 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _529__204
timestamp 1666464484
transform 1 0 25760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _529_
timestamp 1666464484
transform 1 0 27324 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _530_
timestamp 1666464484
transform 1 0 27600 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _530__205
timestamp 1666464484
transform 1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _531_
timestamp 1666464484
transform 1 0 29716 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _531__206
timestamp 1666464484
transform 1 0 25116 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _532_
timestamp 1666464484
transform 1 0 29164 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _532__207
timestamp 1666464484
transform 1 0 28980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _533_
timestamp 1666464484
transform 1 0 29348 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _533__208
timestamp 1666464484
transform 1 0 28704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _534__209
timestamp 1666464484
transform 1 0 28520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _534_
timestamp 1666464484
transform 1 0 29440 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _535__210
timestamp 1666464484
transform 1 0 29808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _535_
timestamp 1666464484
transform 1 0 29900 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _536__211
timestamp 1666464484
transform 1 0 25944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _536_
timestamp 1666464484
transform 1 0 29900 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _537_
timestamp 1666464484
transform 1 0 29900 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _537__212
timestamp 1666464484
transform 1 0 26404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _538__213
timestamp 1666464484
transform -1 0 30728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _538_
timestamp 1666464484
transform 1 0 30452 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _539_
timestamp 1666464484
transform 1 0 30912 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _539__214
timestamp 1666464484
transform -1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _540__215
timestamp 1666464484
transform -1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _540_
timestamp 1666464484
transform -1 0 34224 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _541__216
timestamp 1666464484
transform -1 0 34132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _541_
timestamp 1666464484
transform -1 0 33488 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _542__217
timestamp 1666464484
transform 1 0 32292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _542_
timestamp 1666464484
transform -1 0 34224 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _543__218
timestamp 1666464484
transform -1 0 35144 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _543_
timestamp 1666464484
transform -1 0 34132 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _544__219
timestamp 1666464484
transform -1 0 35788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _544_
timestamp 1666464484
transform -1 0 34592 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _545__220
timestamp 1666464484
transform -1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _545_
timestamp 1666464484
transform -1 0 34408 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _546__221
timestamp 1666464484
transform -1 0 37076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _546_
timestamp 1666464484
transform -1 0 36800 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _547__222
timestamp 1666464484
transform 1 0 33580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _547_
timestamp 1666464484
transform -1 0 35420 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _548_
timestamp 1666464484
transform -1 0 36524 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _548__223
timestamp 1666464484
transform 1 0 36156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _549__224
timestamp 1666464484
transform -1 0 37720 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _549_
timestamp 1666464484
transform -1 0 36524 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _550_
timestamp 1666464484
transform 1 0 34132 0 -1 52224
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _550__225
timestamp 1666464484
transform -1 0 34408 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 3956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1666464484
transform -1 0 28060 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1666464484
transform -1 0 30452 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 32292 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1666464484
transform 1 0 34408 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1666464484
transform -1 0 31832 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1666464484
transform 1 0 35972 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1666464484
transform 1 0 37444 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1666464484
transform 1 0 40020 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1666464484
transform -1 0 40572 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1666464484
transform 1 0 45816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1666464484
transform -1 0 43792 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1666464484
transform 1 0 44252 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1666464484
transform -1 0 46000 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1666464484
transform 1 0 47748 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1666464484
transform 1 0 48392 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1666464484
transform 1 0 50324 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 51612 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1666464484
transform 1 0 52900 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1666464484
transform -1 0 54280 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1666464484
transform -1 0 55844 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_37
timestamp 1666464484
transform -1 0 50600 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_38
timestamp 1666464484
transform -1 0 51888 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_39
timestamp 1666464484
transform -1 0 53268 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_40
timestamp 1666464484
transform -1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_41
timestamp 1666464484
transform -1 0 56488 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_42
timestamp 1666464484
transform -1 0 6808 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_43
timestamp 1666464484
transform -1 0 8004 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_44
timestamp 1666464484
transform -1 0 9568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_45
timestamp 1666464484
transform -1 0 30268 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_46
timestamp 1666464484
transform 1 0 31096 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_47
timestamp 1666464484
transform -1 0 34040 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_48
timestamp 1666464484
transform -1 0 35144 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_49
timestamp 1666464484
transform -1 0 36340 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_50
timestamp 1666464484
transform -1 0 37720 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_51
timestamp 1666464484
transform -1 0 41124 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_52
timestamp 1666464484
transform -1 0 39928 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_53
timestamp 1666464484
transform -1 0 45448 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_54
timestamp 1666464484
transform -1 0 43884 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_55
timestamp 1666464484
transform -1 0 47288 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_56
timestamp 1666464484
transform -1 0 47380 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_57
timestamp 1666464484
transform -1 0 47288 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_58
timestamp 1666464484
transform -1 0 48208 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_59
timestamp 1666464484
transform -1 0 49772 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_60
timestamp 1666464484
transform -1 0 51244 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_61
timestamp 1666464484
transform -1 0 52532 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_62
timestamp 1666464484
transform -1 0 53912 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_63
timestamp 1666464484
transform -1 0 55752 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_64
timestamp 1666464484
transform -1 0 57132 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_65
timestamp 1666464484
transform -1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_66
timestamp 1666464484
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_67
timestamp 1666464484
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_68
timestamp 1666464484
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_69
timestamp 1666464484
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_70
timestamp 1666464484
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_71
timestamp 1666464484
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_72
timestamp 1666464484
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_73
timestamp 1666464484
transform -1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_74
timestamp 1666464484
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_75
timestamp 1666464484
transform 1 0 18676 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_76
timestamp 1666464484
transform -1 0 20700 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_77
timestamp 1666464484
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_78
timestamp 1666464484
transform 1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_79
timestamp 1666464484
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_80
timestamp 1666464484
transform -1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_81
timestamp 1666464484
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_82
timestamp 1666464484
transform 1 0 21252 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_83
timestamp 1666464484
transform -1 0 22632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_84
timestamp 1666464484
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_85
timestamp 1666464484
transform 1 0 21252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_86
timestamp 1666464484
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_87
timestamp 1666464484
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_88
timestamp 1666464484
transform -1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_89
timestamp 1666464484
transform 1 0 23184 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_90
timestamp 1666464484
transform 1 0 20608 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_91
timestamp 1666464484
transform 1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_92
timestamp 1666464484
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_93
timestamp 1666464484
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_94
timestamp 1666464484
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_95
timestamp 1666464484
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_96
timestamp 1666464484
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_97
timestamp 1666464484
transform -1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_98
timestamp 1666464484
transform -1 0 39008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_99
timestamp 1666464484
transform -1 0 38088 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_100
timestamp 1666464484
transform -1 0 37720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_101
timestamp 1666464484
transform -1 0 39008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_102
timestamp 1666464484
transform -1 0 40296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_103
timestamp 1666464484
transform -1 0 38732 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_104
timestamp 1666464484
transform -1 0 39652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_105
timestamp 1666464484
transform -1 0 38364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_106
timestamp 1666464484
transform -1 0 39376 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_107
timestamp 1666464484
transform -1 0 40296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_108
timestamp 1666464484
transform -1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_109
timestamp 1666464484
transform -1 0 39008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_110
timestamp 1666464484
transform -1 0 41584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_111
timestamp 1666464484
transform -1 0 40940 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_112
timestamp 1666464484
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_113
timestamp 1666464484
transform -1 0 39744 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_114
timestamp 1666464484
transform -1 0 41584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_115
timestamp 1666464484
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_116
timestamp 1666464484
transform -1 0 42872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_117
timestamp 1666464484
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_118
timestamp 1666464484
transform -1 0 42872 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_119
timestamp 1666464484
transform -1 0 42228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_120
timestamp 1666464484
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_121
timestamp 1666464484
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_122
timestamp 1666464484
transform -1 0 42872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_123
timestamp 1666464484
transform -1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_124
timestamp 1666464484
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_125
timestamp 1666464484
transform -1 0 44160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_126
timestamp 1666464484
transform -1 0 44160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_127
timestamp 1666464484
transform -1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_128
timestamp 1666464484
transform -1 0 45448 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_129
timestamp 1666464484
transform -1 0 45448 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_130
timestamp 1666464484
transform -1 0 46092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_131
timestamp 1666464484
transform -1 0 45448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_132
timestamp 1666464484
transform -1 0 46736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_133
timestamp 1666464484
transform -1 0 46092 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_134
timestamp 1666464484
transform -1 0 46092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_135
timestamp 1666464484
transform -1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_136
timestamp 1666464484
transform -1 0 46736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_137
timestamp 1666464484
transform -1 0 48024 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_138
timestamp 1666464484
transform -1 0 47380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_139
timestamp 1666464484
transform -1 0 48668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_140
timestamp 1666464484
transform -1 0 48024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_141
timestamp 1666464484
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_142
timestamp 1666464484
transform -1 0 49312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_143
timestamp 1666464484
transform -1 0 48668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_144
timestamp 1666464484
transform -1 0 48668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_145
timestamp 1666464484
transform -1 0 49312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_146
timestamp 1666464484
transform -1 0 50600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_147
timestamp 1666464484
transform -1 0 49956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_148
timestamp 1666464484
transform -1 0 49404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_149
timestamp 1666464484
transform -1 0 51244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_150
timestamp 1666464484
transform -1 0 50600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_151
timestamp 1666464484
transform -1 0 51888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_152
timestamp 1666464484
transform -1 0 51244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_153
timestamp 1666464484
transform -1 0 50784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_154
timestamp 1666464484
transform -1 0 51888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_155
timestamp 1666464484
transform -1 0 51428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_156
timestamp 1666464484
transform -1 0 53176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_157
timestamp 1666464484
transform -1 0 52072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_158
timestamp 1666464484
transform -1 0 53820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_159
timestamp 1666464484
transform -1 0 53176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_160
timestamp 1666464484
transform -1 0 54464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_161
timestamp 1666464484
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_162
timestamp 1666464484
transform -1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_163
timestamp 1666464484
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_164
timestamp 1666464484
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_165
timestamp 1666464484
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_166
timestamp 1666464484
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_167
timestamp 1666464484
transform -1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_168
timestamp 1666464484
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_169
timestamp 1666464484
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_170
timestamp 1666464484
transform -1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_171
timestamp 1666464484
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_172
timestamp 1666464484
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_173
timestamp 1666464484
transform -1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_174
timestamp 1666464484
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_175
timestamp 1666464484
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_176
timestamp 1666464484
transform -1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_177
timestamp 1666464484
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_178
timestamp 1666464484
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_179
timestamp 1666464484
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_180
timestamp 1666464484
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_181
timestamp 1666464484
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_182
timestamp 1666464484
transform -1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_183
timestamp 1666464484
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_184
timestamp 1666464484
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_185
timestamp 1666464484
transform -1 0 15272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_186
timestamp 1666464484
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_187
timestamp 1666464484
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_188
timestamp 1666464484
transform -1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_189
timestamp 1666464484
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_190
timestamp 1666464484
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_191
timestamp 1666464484
transform -1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_192
timestamp 1666464484
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_193
timestamp 1666464484
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_226
timestamp 1666464484
transform -1 0 4968 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_227
timestamp 1666464484
transform -1 0 6164 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_228
timestamp 1666464484
transform 1 0 7084 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_229
timestamp 1666464484
transform 1 0 8372 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_230
timestamp 1666464484
transform -1 0 10304 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_231
timestamp 1666464484
transform -1 0 11868 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_232
timestamp 1666464484
transform -1 0 13064 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_233
timestamp 1666464484
transform -1 0 14628 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_234
timestamp 1666464484
transform -1 0 16008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_235
timestamp 1666464484
transform -1 0 17388 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_236
timestamp 1666464484
transform -1 0 18768 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_237
timestamp 1666464484
transform -1 0 20148 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_238
timestamp 1666464484
transform -1 0 21344 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_239
timestamp 1666464484
transform -1 0 22908 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_240
timestamp 1666464484
transform 1 0 21252 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_241
timestamp 1666464484
transform 1 0 22724 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_242
timestamp 1666464484
transform 1 0 26312 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_243
timestamp 1666464484
transform 1 0 27692 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_244
timestamp 1666464484
transform 1 0 28428 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_245
timestamp 1666464484
transform -1 0 31096 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_246
timestamp 1666464484
transform -1 0 33396 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_247
timestamp 1666464484
transform -1 0 36156 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_248
timestamp 1666464484
transform -1 0 39008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_249
timestamp 1666464484
transform -1 0 36984 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_250
timestamp 1666464484
transform -1 0 42412 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_251
timestamp 1666464484
transform -1 0 40296 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_252
timestamp 1666464484
transform -1 0 43700 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_253
timestamp 1666464484
transform -1 0 46644 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_254
timestamp 1666464484
transform -1 0 46736 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_255
timestamp 1666464484
transform -1 0 46644 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_256
timestamp 1666464484
transform -1 0 48024 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_257
timestamp 1666464484
transform -1 0 49312 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  macro_nodecap_258
timestamp 1666464484
transform -1 0 49128 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1666464484
transform -1 0 5520 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1666464484
transform -1 0 19780 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1666464484
transform -1 0 20700 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1666464484
transform -1 0 22080 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1666464484
transform -1 0 22540 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1666464484
transform -1 0 23276 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1666464484
transform 1 0 25852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1666464484
transform 1 0 27232 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1666464484
transform -1 0 28980 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1666464484
transform -1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1666464484
transform -1 0 12420 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1666464484
transform -1 0 13800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1666464484
transform -1 0 15180 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1666464484
transform -1 0 17204 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1666464484
transform -1 0 17940 0 -1 57664
box -38 -48 406 592
<< labels >>
flabel metal2 s 3698 59200 3754 60000 0 FreeSans 224 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 4158 59200 4214 60000 0 FreeSans 224 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 17958 59200 18014 60000 0 FreeSans 224 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 19338 59200 19394 60000 0 FreeSans 224 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 20718 59200 20774 60000 0 FreeSans 224 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 23478 59200 23534 60000 0 FreeSans 224 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 24858 59200 24914 60000 0 FreeSans 224 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 26238 59200 26294 60000 0 FreeSans 224 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 27618 59200 27674 60000 0 FreeSans 224 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 28998 59200 29054 60000 0 FreeSans 224 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 30378 59200 30434 60000 0 FreeSans 224 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 5538 59200 5594 60000 0 FreeSans 224 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 31758 59200 31814 60000 0 FreeSans 224 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 33138 59200 33194 60000 0 FreeSans 224 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 34518 59200 34574 60000 0 FreeSans 224 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 35898 59200 35954 60000 0 FreeSans 224 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 37278 59200 37334 60000 0 FreeSans 224 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 38658 59200 38714 60000 0 FreeSans 224 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 40038 59200 40094 60000 0 FreeSans 224 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 41418 59200 41474 60000 0 FreeSans 224 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 42798 59200 42854 60000 0 FreeSans 224 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 44178 59200 44234 60000 0 FreeSans 224 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6918 59200 6974 60000 0 FreeSans 224 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 46938 59200 46994 60000 0 FreeSans 224 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 48318 59200 48374 60000 0 FreeSans 224 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 49698 59200 49754 60000 0 FreeSans 224 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 51078 59200 51134 60000 0 FreeSans 224 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 52458 59200 52514 60000 0 FreeSans 224 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 53838 59200 53894 60000 0 FreeSans 224 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 55218 59200 55274 60000 0 FreeSans 224 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 8298 59200 8354 60000 0 FreeSans 224 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 9678 59200 9734 60000 0 FreeSans 224 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 11058 59200 11114 60000 0 FreeSans 224 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 12438 59200 12494 60000 0 FreeSans 224 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 13818 59200 13874 60000 0 FreeSans 224 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 15198 59200 15254 60000 0 FreeSans 224 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 16578 59200 16634 60000 0 FreeSans 224 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 4618 59200 4674 60000 0 FreeSans 224 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 18418 59200 18474 60000 0 FreeSans 224 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 19798 59200 19854 60000 0 FreeSans 224 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 21178 59200 21234 60000 0 FreeSans 224 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 22558 59200 22614 60000 0 FreeSans 224 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 23938 59200 23994 60000 0 FreeSans 224 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 25318 59200 25374 60000 0 FreeSans 224 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 26698 59200 26754 60000 0 FreeSans 224 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 28078 59200 28134 60000 0 FreeSans 224 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 29458 59200 29514 60000 0 FreeSans 224 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 30838 59200 30894 60000 0 FreeSans 224 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 5998 59200 6054 60000 0 FreeSans 224 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 32218 59200 32274 60000 0 FreeSans 224 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 33598 59200 33654 60000 0 FreeSans 224 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 34978 59200 35034 60000 0 FreeSans 224 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 36358 59200 36414 60000 0 FreeSans 224 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 39118 59200 39174 60000 0 FreeSans 224 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 40498 59200 40554 60000 0 FreeSans 224 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 41878 59200 41934 60000 0 FreeSans 224 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 43258 59200 43314 60000 0 FreeSans 224 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 44638 59200 44694 60000 0 FreeSans 224 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 7378 59200 7434 60000 0 FreeSans 224 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 46018 59200 46074 60000 0 FreeSans 224 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 47398 59200 47454 60000 0 FreeSans 224 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 48778 59200 48834 60000 0 FreeSans 224 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 50158 59200 50214 60000 0 FreeSans 224 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 51538 59200 51594 60000 0 FreeSans 224 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 52918 59200 52974 60000 0 FreeSans 224 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 54298 59200 54354 60000 0 FreeSans 224 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 55678 59200 55734 60000 0 FreeSans 224 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8758 59200 8814 60000 0 FreeSans 224 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 10138 59200 10194 60000 0 FreeSans 224 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 11518 59200 11574 60000 0 FreeSans 224 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 12898 59200 12954 60000 0 FreeSans 224 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 15658 59200 15714 60000 0 FreeSans 224 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 17038 59200 17094 60000 0 FreeSans 224 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 5078 59200 5134 60000 0 FreeSans 224 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 18878 59200 18934 60000 0 FreeSans 224 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 20258 59200 20314 60000 0 FreeSans 224 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 21638 59200 21694 60000 0 FreeSans 224 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 23018 59200 23074 60000 0 FreeSans 224 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 24398 59200 24454 60000 0 FreeSans 224 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 25778 59200 25834 60000 0 FreeSans 224 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 27158 59200 27214 60000 0 FreeSans 224 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 28538 59200 28594 60000 0 FreeSans 224 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 31298 59200 31354 60000 0 FreeSans 224 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 32678 59200 32734 60000 0 FreeSans 224 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 34058 59200 34114 60000 0 FreeSans 224 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 35438 59200 35494 60000 0 FreeSans 224 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 36818 59200 36874 60000 0 FreeSans 224 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 38198 59200 38254 60000 0 FreeSans 224 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 39578 59200 39634 60000 0 FreeSans 224 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 40958 59200 41014 60000 0 FreeSans 224 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 42338 59200 42394 60000 0 FreeSans 224 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 43718 59200 43774 60000 0 FreeSans 224 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 45098 59200 45154 60000 0 FreeSans 224 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7838 59200 7894 60000 0 FreeSans 224 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 46478 59200 46534 60000 0 FreeSans 224 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 47858 59200 47914 60000 0 FreeSans 224 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 49238 59200 49294 60000 0 FreeSans 224 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 50618 59200 50674 60000 0 FreeSans 224 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 51998 59200 52054 60000 0 FreeSans 224 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 54758 59200 54814 60000 0 FreeSans 224 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 56138 59200 56194 60000 0 FreeSans 224 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 9218 59200 9274 60000 0 FreeSans 224 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 10598 59200 10654 60000 0 FreeSans 224 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 11978 59200 12034 60000 0 FreeSans 224 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 13358 59200 13414 60000 0 FreeSans 224 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 14738 59200 14794 60000 0 FreeSans 224 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 16118 59200 16174 60000 0 FreeSans 224 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 17498 59200 17554 60000 0 FreeSans 224 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 115 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 116 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 117 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 118 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 119 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 120 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 121 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 122 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 123 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 124 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 125 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 126 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 127 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 128 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 129 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 130 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 131 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 132 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 133 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 134 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 135 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 136 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 137 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 138 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 139 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 140 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 141 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 142 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 143 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 144 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 145 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 146 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 147 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 148 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 149 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 150 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 151 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 152 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 153 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 154 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 155 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 156 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 157 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 158 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 159 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 160 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 161 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 162 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 163 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 164 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 165 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 166 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 167 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 168 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 169 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 170 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 171 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 172 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 173 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 174 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 175 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 176 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 177 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 178 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 179 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 180 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 181 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 182 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 183 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 184 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 185 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 186 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 187 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 188 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 189 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 191 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 192 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 193 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 194 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 195 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 196 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 197 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 198 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 199 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 200 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 201 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 202 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 203 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 204 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 205 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 206 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 207 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 208 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 209 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 210 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 211 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 212 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 213 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 214 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 215 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 216 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 217 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 218 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 219 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 220 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 221 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 222 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 223 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 224 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 225 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 226 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 227 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 228 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 229 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 230 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 231 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 232 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 233 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 234 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 235 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 236 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 237 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 238 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 239 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 240 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 241 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 242 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 243 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 244 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 245 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 246 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 247 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 248 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 249 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 250 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 251 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 252 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 253 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 254 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 255 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 256 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 257 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 258 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 259 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 260 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 261 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 262 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 263 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 264 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 265 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 266 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 267 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 268 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 269 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 270 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 271 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 272 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 273 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 274 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 275 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 276 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 277 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 278 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 279 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 280 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 281 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 282 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 283 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 284 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 285 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 286 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 287 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 288 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 289 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 290 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 291 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 292 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 293 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 294 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 295 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 296 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 297 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 298 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 299 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 300 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 301 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 302 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 303 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 304 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 305 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 306 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 307 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 308 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 309 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 310 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 311 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 312 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 313 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 314 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 315 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 316 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 317 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 319 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 320 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 321 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 322 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 323 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 324 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 325 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 326 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 327 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 328 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 329 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 330 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 331 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 332 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 333 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 334 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 335 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 336 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 337 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 338 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 339 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 340 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 341 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 342 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 343 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 344 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 345 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 346 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 347 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 348 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 349 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 350 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 351 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 352 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 353 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 354 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 355 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 356 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 357 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 358 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 359 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 360 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 361 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 362 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 363 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 364 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 365 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 366 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 367 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 368 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 369 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 370 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 371 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 372 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 373 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 374 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 375 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 376 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 377 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 378 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 379 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 380 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 381 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 382 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 383 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 384 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 385 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 386 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 387 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 388 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 389 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 390 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 391 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 392 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 393 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 394 nsew signal input
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 395 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 396 nsew signal input
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 397 nsew signal input
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 398 nsew signal input
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 399 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 400 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 401 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 402 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 403 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 404 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 405 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 406 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 407 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 408 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 409 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 410 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 411 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 412 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 413 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 414 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 415 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 416 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 417 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 418 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 419 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 420 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 421 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 422 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 423 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 424 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 425 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 426 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 427 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 428 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 429 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 430 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 431 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 432 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 433 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 434 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 435 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 436 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 437 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 438 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 439 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 440 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 441 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 442 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 443 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 444 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 445 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 447 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 448 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 449 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 450 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 451 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 452 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 453 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 454 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 455 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 456 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 457 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 458 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 459 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 460 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 461 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 462 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 463 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 464 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 465 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 466 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 467 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 468 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 469 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 470 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 471 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 472 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 473 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 474 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 475 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 476 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 477 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 478 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 479 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 480 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 481 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 482 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 483 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 484 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 485 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 486 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 487 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 488 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 489 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 490 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 491 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 492 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 493 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 494 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 495 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 496 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 497 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 498 nsew signal input
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 499 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 500 nsew ground bidirectional
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wb_clk_i
port 501 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wb_rst_i
port 502 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 503 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 504 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 505 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 506 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 507 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 508 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 509 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 510 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 511 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 512 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 513 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 514 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 515 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 516 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 517 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 518 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 519 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 520 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 521 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 522 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 523 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 524 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 525 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 526 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 527 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 528 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 529 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 530 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 531 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 532 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 533 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 534 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 535 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 536 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 537 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 538 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 539 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 540 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 541 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 542 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 543 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 544 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 545 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 546 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 547 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 548 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 549 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 550 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 551 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 552 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 553 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 554 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 555 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 556 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 557 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 558 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 559 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 560 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 561 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 562 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 563 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 564 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 565 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 566 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 567 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 568 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 569 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 570 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 571 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 572 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 573 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 574 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 575 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 576 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 577 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 578 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 579 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 580 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 581 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 582 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 583 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 584 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 585 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 586 nsew signal tristate
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 587 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 588 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 589 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 590 nsew signal tristate
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 591 nsew signal tristate
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 592 nsew signal tristate
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 593 nsew signal tristate
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 594 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 595 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 596 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 597 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 598 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 599 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 600 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 601 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 602 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 603 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 604 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 605 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_we_i
port 606 nsew signal input
rlabel metal1 29992 57120 29992 57120 0 vccd1
rlabel metal1 29992 57664 29992 57664 0 vssd1
rlabel metal1 35604 55250 35604 55250 0 _000_
rlabel metal1 35144 55386 35144 55386 0 _001_
rlabel via2 30314 55675 30314 55675 0 _002_
rlabel metal1 29348 55794 29348 55794 0 _003_
rlabel metal1 34868 53754 34868 53754 0 _004_
rlabel metal1 34914 53992 34914 53992 0 _005_
rlabel metal1 29348 54298 29348 54298 0 _006_
rlabel metal1 33856 53754 33856 53754 0 _007_
rlabel metal1 33534 53958 33534 53958 0 _008_
rlabel metal1 33028 53754 33028 53754 0 _009_
rlabel metal1 32338 54094 32338 54094 0 _010_
rlabel metal1 32522 54842 32522 54842 0 _011_
rlabel metal2 31142 54196 31142 54196 0 _012_
rlabel metal2 29854 54842 29854 54842 0 _013_
rlabel metal2 29762 54978 29762 54978 0 _014_
rlabel metal1 28934 55726 28934 55726 0 _015_
rlabel metal1 33051 55930 33051 55930 0 _016_
rlabel metal2 28474 56134 28474 56134 0 _017_
rlabel metal1 28888 56338 28888 56338 0 _018_
rlabel metal1 28060 56474 28060 56474 0 _019_
rlabel metal1 44160 55726 44160 55726 0 _020_
rlabel metal1 44804 55726 44804 55726 0 _021_
rlabel metal1 39100 56338 39100 56338 0 _022_
rlabel metal2 39146 56304 39146 56304 0 _023_
rlabel metal2 44206 54502 44206 54502 0 _024_
rlabel metal1 39698 54706 39698 54706 0 _025_
rlabel metal1 38939 55318 38939 55318 0 _026_
rlabel metal2 42734 54672 42734 54672 0 _027_
rlabel metal2 42642 54332 42642 54332 0 _028_
rlabel metal1 42136 54502 42136 54502 0 _029_
rlabel metal2 41262 54400 41262 54400 0 _030_
rlabel metal1 41998 54638 41998 54638 0 _031_
rlabel metal2 40434 55454 40434 55454 0 _032_
rlabel metal1 38456 56270 38456 56270 0 _033_
rlabel metal2 38226 55046 38226 55046 0 _034_
rlabel metal1 38732 55182 38732 55182 0 _035_
rlabel metal1 38410 56780 38410 56780 0 _036_
rlabel metal1 35466 56780 35466 56780 0 _037_
rlabel metal1 36662 56882 36662 56882 0 _038_
rlabel metal1 28336 57018 28336 57018 0 _039_
rlabel metal1 33580 56338 33580 56338 0 _040_
rlabel metal1 33074 56848 33074 56848 0 _041_
rlabel metal2 32338 56508 32338 56508 0 _042_
rlabel metal2 30590 57154 30590 57154 0 _043_
rlabel metal2 36754 57052 36754 57052 0 _044_
rlabel metal2 41078 57222 41078 57222 0 _045_
rlabel metal2 40526 57052 40526 57052 0 _046_
rlabel metal2 40066 56729 40066 56729 0 _047_
rlabel metal2 24058 56474 24058 56474 0 _048_
rlabel metal2 23598 56814 23598 56814 0 _049_
rlabel metal2 32522 54332 32522 54332 0 _050_
rlabel metal1 33074 54298 33074 54298 0 _051_
rlabel metal1 33948 56338 33948 56338 0 _052_
rlabel metal2 33166 55930 33166 55930 0 _053_
rlabel metal1 32752 55862 32752 55862 0 _054_
rlabel metal2 41170 54604 41170 54604 0 _055_
rlabel metal1 41676 54298 41676 54298 0 _056_
rlabel metal1 43102 55930 43102 55930 0 _057_
rlabel metal1 42136 56338 42136 56338 0 _058_
rlabel metal1 25576 55726 25576 55726 0 _059_
rlabel metal1 25116 55726 25116 55726 0 _060_
rlabel metal2 25530 55692 25530 55692 0 _061_
rlabel metal1 31694 55658 31694 55658 0 _062_
rlabel metal2 31418 55556 31418 55556 0 _063_
rlabel metal2 31050 54944 31050 54944 0 _064_
rlabel metal1 31004 55386 31004 55386 0 _065_
rlabel metal2 30958 55284 30958 55284 0 _066_
rlabel metal1 27997 56338 27997 56338 0 _067_
rlabel metal1 42274 56406 42274 56406 0 _068_
rlabel metal2 40526 56134 40526 56134 0 _069_
rlabel metal2 40250 55046 40250 55046 0 _070_
rlabel metal1 40112 55930 40112 55930 0 _071_
rlabel metal1 40115 55386 40115 55386 0 _072_
rlabel via2 40802 56253 40802 56253 0 _073_
rlabel metal2 26634 55760 26634 55760 0 _074_
rlabel metal2 27186 55420 27186 55420 0 _075_
rlabel metal1 28888 54162 28888 54162 0 _076_
rlabel metal2 28566 54298 28566 54298 0 _077_
rlabel metal1 26818 56848 26818 56848 0 _078_
rlabel metal1 28750 56780 28750 56780 0 _079_
rlabel metal1 32775 56746 32775 56746 0 _080_
rlabel metal1 30130 56882 30130 56882 0 _081_
rlabel metal2 28842 57086 28842 57086 0 _082_
rlabel metal1 37444 55726 37444 55726 0 _083_
rlabel metal2 36846 55964 36846 55964 0 _084_
rlabel metal2 36938 56134 36938 56134 0 _085_
rlabel metal2 43378 57052 43378 57052 0 _086_
rlabel metal2 36570 56916 36570 56916 0 _087_
rlabel metal2 36478 56712 36478 56712 0 _088_
rlabel metal1 25208 6766 25208 6766 0 _089_
rlabel metal1 33396 5678 33396 5678 0 _090_
rlabel metal2 25806 3026 25806 3026 0 _091_
rlabel metal1 24702 4692 24702 4692 0 _092_
rlabel metal2 25254 6188 25254 6188 0 _093_
rlabel metal1 24288 4046 24288 4046 0 _094_
rlabel metal1 23138 2550 23138 2550 0 _095_
rlabel metal1 23414 2618 23414 2618 0 _096_
rlabel metal1 25392 4522 25392 4522 0 _097_
rlabel metal2 27370 5950 27370 5950 0 _098_
rlabel metal2 27554 5916 27554 5916 0 _099_
rlabel metal1 27600 6834 27600 6834 0 _100_
rlabel metal2 26082 4216 26082 4216 0 _101_
rlabel metal2 24610 2652 24610 2652 0 _102_
rlabel metal1 25093 3366 25093 3366 0 _103_
rlabel metal1 24426 2618 24426 2618 0 _104_
rlabel metal2 29026 2720 29026 2720 0 _105_
rlabel metal1 29256 7718 29256 7718 0 _106_
rlabel metal2 29578 7582 29578 7582 0 _107_
rlabel metal1 29762 3706 29762 3706 0 _108_
rlabel metal2 30498 4114 30498 4114 0 _109_
rlabel metal1 30130 3978 30130 3978 0 _110_
rlabel metal2 30130 2618 30130 2618 0 _111_
rlabel metal1 30636 8330 30636 8330 0 _112_
rlabel metal1 31188 7718 31188 7718 0 _113_
rlabel metal1 35558 2346 35558 2346 0 _114_
rlabel metal1 34822 2618 34822 2618 0 _115_
rlabel metal2 33994 5406 33994 5406 0 _116_
rlabel metal1 34454 4522 34454 4522 0 _117_
rlabel metal1 34362 4012 34362 4012 0 _118_
rlabel metal1 36156 2074 36156 2074 0 _119_
rlabel metal1 36938 3434 36938 3434 0 _120_
rlabel metal2 35650 6018 35650 6018 0 _121_
rlabel metal2 36294 5406 36294 5406 0 _122_
rlabel metal1 37260 3094 37260 3094 0 _123_
rlabel metal1 27876 54570 27876 54570 0 _124_
rlabel metal1 3588 57562 3588 57562 0 io_active
rlabel metal1 28382 55250 28382 55250 0 io_in[18]
rlabel metal1 30360 57426 30360 57426 0 io_in[19]
rlabel metal1 32200 57358 32200 57358 0 io_in[20]
rlabel metal1 33994 55250 33994 55250 0 io_in[21]
rlabel metal2 34546 58388 34546 58388 0 io_in[22]
rlabel metal1 35972 57426 35972 57426 0 io_in[23]
rlabel metal1 37398 57426 37398 57426 0 io_in[24]
rlabel metal1 39376 57426 39376 57426 0 io_in[25]
rlabel metal2 40342 56695 40342 56695 0 io_in[26]
rlabel metal1 46000 56814 46000 56814 0 io_in[27]
rlabel metal1 43286 57426 43286 57426 0 io_in[28]
rlabel metal1 44344 55250 44344 55250 0 io_in[29]
rlabel metal1 45724 57494 45724 57494 0 io_in[30]
rlabel metal1 47380 57358 47380 57358 0 io_in[31]
rlabel metal1 48392 56882 48392 56882 0 io_in[32]
rlabel metal1 50048 57426 50048 57426 0 io_in[33]
rlabel metal1 51382 57426 51382 57426 0 io_in[34]
rlabel metal1 52762 57494 52762 57494 0 io_in[35]
rlabel metal1 54050 57426 54050 57426 0 io_in[36]
rlabel metal1 55522 57426 55522 57426 0 io_in[37]
rlabel metal1 5198 57562 5198 57562 0 io_out[0]
rlabel metal1 19458 57562 19458 57562 0 io_out[10]
rlabel metal1 20378 57562 20378 57562 0 io_out[11]
rlabel metal1 21758 57018 21758 57018 0 io_out[12]
rlabel metal1 22678 57562 22678 57562 0 io_out[13]
rlabel metal1 23276 57290 23276 57290 0 io_out[14]
rlabel metal1 25944 57562 25944 57562 0 io_out[15]
rlabel metal1 27324 57562 27324 57562 0 io_out[16]
rlabel metal1 28658 57562 28658 57562 0 io_out[17]
rlabel metal1 10718 57562 10718 57562 0 io_out[4]
rlabel metal1 12098 57562 12098 57562 0 io_out[5]
rlabel metal1 13478 57562 13478 57562 0 io_out[6]
rlabel metal1 14858 57562 14858 57562 0 io_out[7]
rlabel metal2 16146 58388 16146 58388 0 io_out[8]
rlabel metal1 17618 57562 17618 57562 0 io_out[9]
rlabel metal2 25990 4335 25990 4335 0 la_data_out[32]
rlabel metal2 26450 2404 26450 2404 0 la_data_out[33]
rlabel metal2 26726 2166 26726 2166 0 la_data_out[34]
rlabel metal2 27002 1860 27002 1860 0 la_data_out[35]
rlabel metal2 27278 1775 27278 1775 0 la_data_out[36]
rlabel metal2 27554 1707 27554 1707 0 la_data_out[37]
rlabel metal2 27830 3254 27830 3254 0 la_data_out[38]
rlabel metal2 28106 3798 28106 3798 0 la_data_out[39]
rlabel metal2 28382 2404 28382 2404 0 la_data_out[40]
rlabel metal2 28658 959 28658 959 0 la_data_out[41]
rlabel metal2 28934 2166 28934 2166 0 la_data_out[42]
rlabel metal2 29210 1860 29210 1860 0 la_data_out[43]
rlabel metal2 29486 1792 29486 1792 0 la_data_out[44]
rlabel metal2 29762 3492 29762 3492 0 la_data_out[45]
rlabel metal2 30038 2098 30038 2098 0 la_data_out[46]
rlabel metal2 30314 1775 30314 1775 0 la_data_out[47]
rlabel metal2 30590 2710 30590 2710 0 la_data_out[48]
rlabel metal2 30866 2404 30866 2404 0 la_data_out[49]
rlabel metal2 31142 1860 31142 1860 0 la_data_out[50]
rlabel metal2 31418 3254 31418 3254 0 la_data_out[51]
rlabel metal2 31694 3798 31694 3798 0 la_data_out[52]
rlabel metal1 32154 2958 32154 2958 0 la_data_out[53]
rlabel metal2 32246 2166 32246 2166 0 la_data_out[54]
rlabel metal2 32522 2948 32522 2948 0 la_data_out[55]
rlabel metal2 32798 1761 32798 1761 0 la_data_out[56]
rlabel metal2 33074 2404 33074 2404 0 la_data_out[57]
rlabel metal2 33350 1622 33350 1622 0 la_data_out[58]
rlabel metal1 34270 3570 34270 3570 0 la_data_out[59]
rlabel metal2 33902 3492 33902 3492 0 la_data_out[60]
rlabel metal1 34454 3706 34454 3706 0 la_data_out[61]
rlabel metal1 34546 2958 34546 2958 0 la_data_out[62]
rlabel metal2 34730 1078 34730 1078 0 la_data_out[63]
rlabel metal2 5474 56814 5474 56814 0 net1
rlabel metal1 40710 54842 40710 54842 0 net10
rlabel metal1 35834 4012 35834 4012 0 net100
rlabel metal1 36846 2890 36846 2890 0 net101
rlabel metal1 38226 3366 38226 3366 0 net102
rlabel metal2 36800 3332 36800 3332 0 net103
rlabel metal1 38180 3162 38180 3162 0 net104
rlabel metal1 37674 3978 37674 3978 0 net105
rlabel metal2 37490 1095 37490 1095 0 net106
rlabel metal1 38640 2890 38640 2890 0 net107
rlabel metal2 38042 1622 38042 1622 0 net108
rlabel metal1 38548 3910 38548 3910 0 net109
rlabel metal1 42872 55726 42872 55726 0 net11
rlabel metal2 38594 1588 38594 1588 0 net110
rlabel metal1 39790 2958 39790 2958 0 net111
rlabel metal1 39606 3638 39606 3638 0 net112
rlabel metal1 39468 3910 39468 3910 0 net113
rlabel metal1 40526 2890 40526 2890 0 net114
rlabel metal1 40342 3570 40342 3570 0 net115
rlabel metal1 42642 2380 42642 2380 0 net116
rlabel metal1 40940 3502 40940 3502 0 net117
rlabel metal2 40802 1860 40802 1860 0 net118
rlabel metal2 41078 2200 41078 2200 0 net119
rlabel metal1 43562 57358 43562 57358 0 net12
rlabel metal2 41446 1955 41446 1955 0 net120
rlabel metal2 41630 1826 41630 1826 0 net121
rlabel metal2 41906 2166 41906 2166 0 net122
rlabel metal2 42182 1656 42182 1656 0 net123
rlabel metal2 42458 2132 42458 2132 0 net124
rlabel metal2 42734 1894 42734 1894 0 net125
rlabel metal2 43010 2166 43010 2166 0 net126
rlabel metal2 43286 1860 43286 1860 0 net127
rlabel metal2 43562 1622 43562 1622 0 net128
rlabel metal2 43838 1792 43838 1792 0 net129
rlabel metal1 39238 55624 39238 55624 0 net13
rlabel metal2 44114 1554 44114 1554 0 net130
rlabel metal2 44390 2132 44390 2132 0 net131
rlabel metal2 44666 1656 44666 1656 0 net132
rlabel metal2 44942 1826 44942 1826 0 net133
rlabel metal2 45218 2200 45218 2200 0 net134
rlabel metal2 45494 1792 45494 1792 0 net135
rlabel metal2 45770 2132 45770 2132 0 net136
rlabel metal2 46046 1588 46046 1588 0 net137
rlabel metal2 46322 2098 46322 2098 0 net138
rlabel metal2 46598 1622 46598 1622 0 net139
rlabel metal1 41101 54638 41101 54638 0 net14
rlabel metal2 46874 1792 46874 1792 0 net140
rlabel metal2 47150 2200 47150 2200 0 net141
rlabel metal2 47426 1554 47426 1554 0 net142
rlabel metal2 47702 1826 47702 1826 0 net143
rlabel metal2 47978 2132 47978 2132 0 net144
rlabel metal2 48254 1792 48254 1792 0 net145
rlabel metal2 48530 1656 48530 1656 0 net146
rlabel metal2 48806 1860 48806 1860 0 net147
rlabel metal2 49082 2132 49082 2132 0 net148
rlabel metal2 49358 1622 49358 1622 0 net149
rlabel metal1 45632 55862 45632 55862 0 net15
rlabel metal2 49634 1826 49634 1826 0 net150
rlabel metal2 49910 1588 49910 1588 0 net151
rlabel metal2 50186 1792 50186 1792 0 net152
rlabel metal2 50462 1299 50462 1299 0 net153
rlabel metal2 50738 1826 50738 1826 0 net154
rlabel metal2 51014 2132 51014 2132 0 net155
rlabel metal2 51290 1554 51290 1554 0 net156
rlabel metal2 51566 2132 51566 2132 0 net157
rlabel metal2 51842 1656 51842 1656 0 net158
rlabel metal2 52118 1792 52118 1792 0 net159
rlabel metal2 45402 56236 45402 56236 0 net16
rlabel metal2 52394 1622 52394 1622 0 net160
rlabel metal2 7682 1588 7682 1588 0 net161
rlabel metal2 8234 1792 8234 1792 0 net162
rlabel metal2 8602 1656 8602 1656 0 net163
rlabel metal2 8970 2132 8970 2132 0 net164
rlabel metal2 9338 1588 9338 1588 0 net165
rlabel metal2 9706 1792 9706 1792 0 net166
rlabel metal2 9982 2132 9982 2132 0 net167
rlabel metal2 10258 1792 10258 1792 0 net168
rlabel metal2 10534 1656 10534 1656 0 net169
rlabel metal1 45310 57426 45310 57426 0 net17
rlabel metal2 10810 2132 10810 2132 0 net170
rlabel metal2 11086 1792 11086 1792 0 net171
rlabel metal2 11362 1792 11362 1792 0 net172
rlabel metal2 11638 2132 11638 2132 0 net173
rlabel metal2 11914 1554 11914 1554 0 net174
rlabel metal2 12190 1588 12190 1588 0 net175
rlabel metal2 12466 2132 12466 2132 0 net176
rlabel metal2 12742 1792 12742 1792 0 net177
rlabel metal2 13018 1588 13018 1588 0 net178
rlabel metal2 13294 2132 13294 2132 0 net179
rlabel metal2 51842 56508 51842 56508 0 net18
rlabel metal2 13570 1792 13570 1792 0 net180
rlabel metal2 13846 1622 13846 1622 0 net181
rlabel metal2 14122 2132 14122 2132 0 net182
rlabel metal2 14398 1860 14398 1860 0 net183
rlabel metal2 14674 1792 14674 1792 0 net184
rlabel metal2 14950 2132 14950 2132 0 net185
rlabel metal2 15226 1656 15226 1656 0 net186
rlabel metal2 15502 1792 15502 1792 0 net187
rlabel metal2 15778 2132 15778 2132 0 net188
rlabel metal2 16054 1588 16054 1588 0 net189
rlabel metal2 53130 56202 53130 56202 0 net19
rlabel metal2 16330 1860 16330 1860 0 net190
rlabel metal2 16606 2132 16606 2132 0 net191
rlabel metal2 16882 1792 16882 1792 0 net192
rlabel metal2 17158 1656 17158 1656 0 net193
rlabel metal2 25070 5916 25070 5916 0 net194
rlabel metal1 24748 4114 24748 4114 0 net195
rlabel metal1 22402 3060 22402 3060 0 net196
rlabel metal2 24794 3230 24794 3230 0 net197
rlabel metal2 25346 4828 25346 4828 0 net198
rlabel metal1 26910 5134 26910 5134 0 net199
rlabel metal2 31970 56814 31970 56814 0 net2
rlabel via1 45785 56338 45785 56338 0 net20
rlabel metal1 27692 5814 27692 5814 0 net200
rlabel metal2 27370 7004 27370 7004 0 net201
rlabel metal2 26910 4420 26910 4420 0 net202
rlabel metal2 25898 3162 25898 3162 0 net203
rlabel metal2 27370 4284 27370 4284 0 net204
rlabel metal1 27646 2924 27646 2924 0 net205
rlabel metal1 25783 2550 25783 2550 0 net206
rlabel metal2 29210 5508 29210 5508 0 net207
rlabel metal1 29164 7310 29164 7310 0 net208
rlabel metal2 29486 5644 29486 5644 0 net209
rlabel metal2 54142 57664 54142 57664 0 net21
rlabel metal2 29946 5168 29946 5168 0 net210
rlabel metal2 26174 4420 26174 4420 0 net211
rlabel metal1 26634 2380 26634 2380 0 net212
rlabel metal2 30498 6800 30498 6800 0 net213
rlabel metal1 31234 6290 31234 6290 0 net214
rlabel metal1 35144 2550 35144 2550 0 net215
rlabel metal1 33672 3502 33672 3502 0 net216
rlabel metal2 34178 5644 34178 5644 0 net217
rlabel metal1 34316 4658 34316 4658 0 net218
rlabel metal1 35052 4046 35052 4046 0 net219
rlabel metal1 6072 57358 6072 57358 0 net22
rlabel metal1 34914 2482 34914 2482 0 net220
rlabel viali 36754 3578 36754 3578 0 net221
rlabel metal2 35374 6528 35374 6528 0 net222
rlabel metal1 36432 4794 36432 4794 0 net223
rlabel metal1 36984 2958 36984 2958 0 net224
rlabel metal2 34178 51748 34178 51748 0 net225
rlabel metal1 4692 57018 4692 57018 0 net226
rlabel metal1 5980 57018 5980 57018 0 net227
rlabel metal1 7360 57426 7360 57426 0 net228
rlabel metal1 8694 57426 8694 57426 0 net229
rlabel metal1 19734 57392 19734 57392 0 net23
rlabel metal1 10120 57426 10120 57426 0 net230
rlabel metal1 11592 57018 11592 57018 0 net231
rlabel metal1 12880 57426 12880 57426 0 net232
rlabel metal1 14352 57018 14352 57018 0 net233
rlabel metal1 15732 57426 15732 57426 0 net234
rlabel metal1 17112 57018 17112 57018 0 net235
rlabel metal1 18492 57426 18492 57426 0 net236
rlabel metal1 19964 57018 19964 57018 0 net237
rlabel metal1 21160 57018 21160 57018 0 net238
rlabel metal1 22632 56338 22632 56338 0 net239
rlabel metal1 20654 57460 20654 57460 0 net24
rlabel metal2 22862 57494 22862 57494 0 net240
rlabel metal1 23552 56950 23552 56950 0 net241
rlabel metal1 26634 54842 26634 54842 0 net242
rlabel metal1 28014 54842 28014 54842 0 net243
rlabel metal1 29072 55182 29072 55182 0 net244
rlabel metal2 30866 58320 30866 58320 0 net245
rlabel metal1 32706 55114 32706 55114 0 net246
rlabel metal1 35190 55930 35190 55930 0 net247
rlabel metal2 38778 56848 38778 56848 0 net248
rlabel metal1 36570 55182 36570 55182 0 net249
rlabel metal2 27186 56372 27186 56372 0 net25
rlabel metal1 39146 56440 39146 56440 0 net250
rlabel metal2 40066 55029 40066 55029 0 net251
rlabel metal2 40572 57324 40572 57324 0 net252
rlabel metal2 46414 56729 46414 56729 0 net253
rlabel metal1 45678 56882 45678 56882 0 net254
rlabel metal1 45540 56202 45540 56202 0 net255
rlabel metal1 46920 57018 46920 57018 0 net256
rlabel metal1 48254 57426 48254 57426 0 net257
rlabel metal1 48852 56338 48852 56338 0 net258
rlabel metal2 33994 57358 33994 57358 0 net26
rlabel metal1 23368 57018 23368 57018 0 net27
rlabel metal2 25162 56100 25162 56100 0 net28
rlabel metal2 27278 56882 27278 56882 0 net29
rlabel metal2 34362 56848 34362 56848 0 net3
rlabel metal1 29394 56882 29394 56882 0 net30
rlabel metal2 21390 57426 21390 57426 0 net31
rlabel via2 12374 57443 12374 57443 0 net32
rlabel metal1 13754 57358 13754 57358 0 net33
rlabel metal1 20562 57528 20562 57528 0 net34
rlabel metal2 17158 56814 17158 56814 0 net35
rlabel metal2 17894 57630 17894 57630 0 net36
rlabel metal1 50278 57018 50278 57018 0 net37
rlabel metal1 51612 57018 51612 57018 0 net38
rlabel metal1 52992 57018 52992 57018 0 net39
rlabel metal2 32706 54740 32706 54740 0 net4
rlabel metal1 54510 57426 54510 57426 0 net40
rlabel metal1 55982 57358 55982 57358 0 net41
rlabel metal1 6532 57018 6532 57018 0 net42
rlabel metal1 7820 57426 7820 57426 0 net43
rlabel metal1 9292 57426 9292 57426 0 net44
rlabel metal1 29992 56338 29992 56338 0 net45
rlabel metal2 31326 58116 31326 58116 0 net46
rlabel metal2 33810 55284 33810 55284 0 net47
rlabel metal1 34868 54842 34868 54842 0 net48
rlabel metal1 36110 55250 36110 55250 0 net49
rlabel metal1 34224 55386 34224 55386 0 net5
rlabel metal1 37490 55216 37490 55216 0 net50
rlabel metal1 39560 55862 39560 55862 0 net51
rlabel metal1 39652 54162 39652 54162 0 net52
rlabel metal2 40986 57793 40986 57793 0 net53
rlabel metal1 43654 55284 43654 55284 0 net54
rlabel metal2 47058 56865 47058 56865 0 net55
rlabel metal1 46138 56950 46138 56950 0 net56
rlabel metal1 46782 56338 46782 56338 0 net57
rlabel metal1 47932 56338 47932 56338 0 net58
rlabel metal1 49404 56338 49404 56338 0 net59
rlabel metal1 34362 54094 34362 54094 0 net6
rlabel metal1 50830 57018 50830 57018 0 net60
rlabel metal1 52164 57018 52164 57018 0 net61
rlabel metal1 53544 57018 53544 57018 0 net62
rlabel metal2 55522 56644 55522 56644 0 net63
rlabel metal1 56534 57426 56534 57426 0 net64
rlabel metal2 17342 2336 17342 2336 0 net65
rlabel metal2 17618 2132 17618 2132 0 net66
rlabel metal2 17894 1622 17894 1622 0 net67
rlabel metal2 18170 1792 18170 1792 0 net68
rlabel metal2 18446 2132 18446 2132 0 net69
rlabel metal1 34638 56372 34638 56372 0 net7
rlabel metal2 18722 1792 18722 1792 0 net70
rlabel metal2 18998 1656 18998 1656 0 net71
rlabel metal2 19274 2132 19274 2132 0 net72
rlabel metal2 19550 1367 19550 1367 0 net73
rlabel metal2 19826 1027 19826 1027 0 net74
rlabel metal2 20102 1826 20102 1826 0 net75
rlabel metal2 20378 2336 20378 2336 0 net76
rlabel metal2 20654 2132 20654 2132 0 net77
rlabel metal2 20930 1860 20930 1860 0 net78
rlabel metal2 21206 1554 21206 1554 0 net79
rlabel metal1 35282 55318 35282 55318 0 net8
rlabel metal2 21482 2676 21482 2676 0 net80
rlabel metal2 21758 2166 21758 2166 0 net81
rlabel metal2 22034 2336 22034 2336 0 net82
rlabel metal2 22310 2676 22310 2676 0 net83
rlabel metal2 22586 1826 22586 1826 0 net84
rlabel metal2 22862 2200 22862 2200 0 net85
rlabel metal2 23138 2370 23138 2370 0 net86
rlabel metal2 23414 1622 23414 1622 0 net87
rlabel metal2 23690 2880 23690 2880 0 net88
rlabel metal2 23966 1571 23966 1571 0 net89
rlabel metal1 40342 57460 40342 57460 0 net9
rlabel metal2 24242 1112 24242 1112 0 net90
rlabel metal2 24518 2234 24518 2234 0 net91
rlabel metal2 24794 1843 24794 1843 0 net92
rlabel metal2 25070 1520 25070 1520 0 net93
rlabel metal2 25346 2370 25346 2370 0 net94
rlabel metal2 25622 1554 25622 1554 0 net95
rlabel metal2 25898 1299 25898 1299 0 net96
rlabel metal2 35006 1520 35006 1520 0 net97
rlabel metal2 35282 1095 35282 1095 0 net98
rlabel metal1 36708 3706 36708 3706 0 net99
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
